-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 29 2019 01:19:43

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "corePackage" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of corePackage
entity corePackage is
port (
    o_UART_TX : out std_logic;
    i_UART_RX : in std_logic;
    i_Clk : in std_logic);
end corePackage;

-- Architecture of corePackage
-- View name is \INTERFACE\
architecture \INTERFACE\ of corePackage is

signal \N__1159\ : std_logic;
signal \N__1158\ : std_logic;
signal \N__1157\ : std_logic;
signal \N__1148\ : std_logic;
signal \N__1147\ : std_logic;
signal \N__1146\ : std_logic;
signal \N__1129\ : std_logic;
signal \N__1126\ : std_logic;
signal \N__1123\ : std_logic;
signal \N__1122\ : std_logic;
signal \N__1121\ : std_logic;
signal \N__1116\ : std_logic;
signal \N__1113\ : std_logic;
signal \N__1108\ : std_logic;
signal \N__1105\ : std_logic;
signal \N__1104\ : std_logic;
signal \N__1099\ : std_logic;
signal \N__1096\ : std_logic;
signal \N__1093\ : std_logic;
signal \N__1092\ : std_logic;
signal \N__1091\ : std_logic;
signal \N__1090\ : std_logic;
signal \N__1089\ : std_logic;
signal \N__1088\ : std_logic;
signal \N__1087\ : std_logic;
signal \N__1084\ : std_logic;
signal \N__1081\ : std_logic;
signal \N__1074\ : std_logic;
signal \N__1071\ : std_logic;
signal \N__1068\ : std_logic;
signal \N__1057\ : std_logic;
signal \N__1054\ : std_logic;
signal \N__1053\ : std_logic;
signal \N__1052\ : std_logic;
signal \N__1051\ : std_logic;
signal \N__1048\ : std_logic;
signal \N__1045\ : std_logic;
signal \N__1042\ : std_logic;
signal \N__1039\ : std_logic;
signal \N__1036\ : std_logic;
signal \N__1027\ : std_logic;
signal \N__1026\ : std_logic;
signal \N__1025\ : std_logic;
signal \N__1024\ : std_logic;
signal \N__1023\ : std_logic;
signal \N__1020\ : std_logic;
signal \N__1019\ : std_logic;
signal \N__1018\ : std_logic;
signal \N__1017\ : std_logic;
signal \N__1014\ : std_logic;
signal \N__1005\ : std_logic;
signal \N__1000\ : std_logic;
signal \N__997\ : std_logic;
signal \N__988\ : std_logic;
signal \N__987\ : std_logic;
signal \N__986\ : std_logic;
signal \N__985\ : std_logic;
signal \N__984\ : std_logic;
signal \N__981\ : std_logic;
signal \N__978\ : std_logic;
signal \N__969\ : std_logic;
signal \N__964\ : std_logic;
signal \N__961\ : std_logic;
signal \N__960\ : std_logic;
signal \N__959\ : std_logic;
signal \N__958\ : std_logic;
signal \N__957\ : std_logic;
signal \N__956\ : std_logic;
signal \N__955\ : std_logic;
signal \N__954\ : std_logic;
signal \N__953\ : std_logic;
signal \N__950\ : std_logic;
signal \N__941\ : std_logic;
signal \N__936\ : std_logic;
signal \N__931\ : std_logic;
signal \N__922\ : std_logic;
signal \N__919\ : std_logic;
signal \N__916\ : std_logic;
signal \N__915\ : std_logic;
signal \N__914\ : std_logic;
signal \N__911\ : std_logic;
signal \N__908\ : std_logic;
signal \N__905\ : std_logic;
signal \N__898\ : std_logic;
signal \N__897\ : std_logic;
signal \N__896\ : std_logic;
signal \N__895\ : std_logic;
signal \N__894\ : std_logic;
signal \N__893\ : std_logic;
signal \N__892\ : std_logic;
signal \N__891\ : std_logic;
signal \N__890\ : std_logic;
signal \N__889\ : std_logic;
signal \N__886\ : std_logic;
signal \N__885\ : std_logic;
signal \N__884\ : std_logic;
signal \N__881\ : std_logic;
signal \N__878\ : std_logic;
signal \N__873\ : std_logic;
signal \N__864\ : std_logic;
signal \N__859\ : std_logic;
signal \N__854\ : std_logic;
signal \N__841\ : std_logic;
signal \N__838\ : std_logic;
signal \N__835\ : std_logic;
signal \N__832\ : std_logic;
signal \N__831\ : std_logic;
signal \N__830\ : std_logic;
signal \N__823\ : std_logic;
signal \N__820\ : std_logic;
signal \N__819\ : std_logic;
signal \N__818\ : std_logic;
signal \N__817\ : std_logic;
signal \N__816\ : std_logic;
signal \N__815\ : std_logic;
signal \N__802\ : std_logic;
signal \N__799\ : std_logic;
signal \N__796\ : std_logic;
signal \N__793\ : std_logic;
signal \N__790\ : std_logic;
signal \N__789\ : std_logic;
signal \N__788\ : std_logic;
signal \N__787\ : std_logic;
signal \N__786\ : std_logic;
signal \N__785\ : std_logic;
signal \N__782\ : std_logic;
signal \N__781\ : std_logic;
signal \N__780\ : std_logic;
signal \N__777\ : std_logic;
signal \N__774\ : std_logic;
signal \N__767\ : std_logic;
signal \N__764\ : std_logic;
signal \N__759\ : std_logic;
signal \N__748\ : std_logic;
signal \N__747\ : std_logic;
signal \N__746\ : std_logic;
signal \N__743\ : std_logic;
signal \N__742\ : std_logic;
signal \N__741\ : std_logic;
signal \N__740\ : std_logic;
signal \N__739\ : std_logic;
signal \N__736\ : std_logic;
signal \N__727\ : std_logic;
signal \N__724\ : std_logic;
signal \N__719\ : std_logic;
signal \N__712\ : std_logic;
signal \N__711\ : std_logic;
signal \N__710\ : std_logic;
signal \N__709\ : std_logic;
signal \N__708\ : std_logic;
signal \N__707\ : std_logic;
signal \N__706\ : std_logic;
signal \N__703\ : std_logic;
signal \N__700\ : std_logic;
signal \N__695\ : std_logic;
signal \N__688\ : std_logic;
signal \N__683\ : std_logic;
signal \N__680\ : std_logic;
signal \N__673\ : std_logic;
signal \N__670\ : std_logic;
signal \N__667\ : std_logic;
signal \N__664\ : std_logic;
signal \N__661\ : std_logic;
signal \N__660\ : std_logic;
signal \N__657\ : std_logic;
signal \N__656\ : std_logic;
signal \N__653\ : std_logic;
signal \N__648\ : std_logic;
signal \N__643\ : std_logic;
signal \N__642\ : std_logic;
signal \N__641\ : std_logic;
signal \N__638\ : std_logic;
signal \N__637\ : std_logic;
signal \N__636\ : std_logic;
signal \N__635\ : std_logic;
signal \N__632\ : std_logic;
signal \N__631\ : std_logic;
signal \N__630\ : std_logic;
signal \N__627\ : std_logic;
signal \N__622\ : std_logic;
signal \N__617\ : std_logic;
signal \N__610\ : std_logic;
signal \N__601\ : std_logic;
signal \N__600\ : std_logic;
signal \N__599\ : std_logic;
signal \N__598\ : std_logic;
signal \N__597\ : std_logic;
signal \N__592\ : std_logic;
signal \N__589\ : std_logic;
signal \N__584\ : std_logic;
signal \N__577\ : std_logic;
signal \N__576\ : std_logic;
signal \N__575\ : std_logic;
signal \N__572\ : std_logic;
signal \N__569\ : std_logic;
signal \N__566\ : std_logic;
signal \N__565\ : std_logic;
signal \N__564\ : std_logic;
signal \N__561\ : std_logic;
signal \N__558\ : std_logic;
signal \N__555\ : std_logic;
signal \N__550\ : std_logic;
signal \N__541\ : std_logic;
signal \N__540\ : std_logic;
signal \N__539\ : std_logic;
signal \N__538\ : std_logic;
signal \N__537\ : std_logic;
signal \N__536\ : std_logic;
signal \N__533\ : std_logic;
signal \N__528\ : std_logic;
signal \N__523\ : std_logic;
signal \N__520\ : std_logic;
signal \N__517\ : std_logic;
signal \N__508\ : std_logic;
signal \N__505\ : std_logic;
signal \N__502\ : std_logic;
signal \N__499\ : std_logic;
signal \N__496\ : std_logic;
signal \N__493\ : std_logic;
signal \N__490\ : std_logic;
signal \N__487\ : std_logic;
signal \N__484\ : std_logic;
signal \N__481\ : std_logic;
signal \N__478\ : std_logic;
signal \N__475\ : std_logic;
signal \N__472\ : std_logic;
signal \N__469\ : std_logic;
signal \N__466\ : std_logic;
signal \N__463\ : std_logic;
signal \N__460\ : std_logic;
signal \N__459\ : std_logic;
signal \N__456\ : std_logic;
signal \N__453\ : std_logic;
signal \N__450\ : std_logic;
signal \N__447\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uartTxInst.N_8_i_cascade_\ : std_logic;
signal \uartTxInst.m11_i_a3_3\ : std_logic;
signal \uartTxInst.m11_i_a3_4\ : std_logic;
signal \uartTxInst.m15_e_5\ : std_logic;
signal \uartTxInst.m15_e_4\ : std_logic;
signal \o_UART_TX_c\ : std_logic;
signal \uartTxInst.un5_rclkcount_ac0_11_cascade_\ : std_logic;
signal \uartTxInst.un5_rclkcount_c4_cascade_\ : std_logic;
signal \uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \uartTxInst.N_17_mux\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_1\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_2\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_5\ : std_logic;
signal \uartTxInst.un2_rclkcount_5_cascade_\ : std_logic;
signal \uartTxInst.rClkCount_RNIOIKC_0Z0Z_3\ : std_logic;
signal \uartTxInst.SUM_N_3_mux_cascade_\ : std_logic;
signal \uartTxInst.un5_rclkcount_c4\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_4\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_3\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_7\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_6\ : std_logic;
signal \uartTxInst.un2_rclkcount_4_cascade_\ : std_logic;
signal \uartTxInst.rTxState_10_0_x2_0_o2_1_0_1_cascade_\ : std_logic;
signal \uartTxInst.un2_rclkcount_5\ : std_logic;
signal \uartTxInst.N_20_cascade_\ : std_logic;
signal \uartTxInst.rBitIndexZ0Z_2\ : std_logic;
signal \uartTxInst.rTxStateZ0Z_1\ : std_logic;
signal \uartTxInst.rTxState_10_0_i_a2_0_1_0_cascade_\ : std_logic;
signal \uartTxInst.SUM_N_3_mux\ : std_logic;
signal \uartTxInst.rTxStateZ0Z_0\ : std_logic;
signal \uartTxInst.rBitIndexZ1Z_0\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_0\ : std_logic;
signal \uartTxInst.rBitIndex_RNO_2Z0Z_1\ : std_logic;
signal \uartTxInst.un2_rclkcount_4\ : std_logic;
signal \uartTxInst.rbitindex15\ : std_logic;
signal \uartTxInst.SUM_i_o2_d_1_cascade_\ : std_logic;
signal \uartTxInst.SUM_i_o2_1_0_1\ : std_logic;
signal \uartTxInst.rBitIndexZ0Z_1\ : std_logic;
signal \i_Clk_c_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \i_Clk_wire\ : std_logic;
signal \o_UART_TX_wire\ : std_logic;

begin
    \i_Clk_wire\ <= i_Clk;
    o_UART_TX <= \o_UART_TX_wire\;

    \i_Clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__1157\,
            GLOBALBUFFEROUTPUT => \i_Clk_c_g\
        );

    \i_Clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1159\,
            DIN => \N__1158\,
            DOUT => \N__1157\,
            PACKAGEPIN => \i_Clk_wire\
        );

    \i_Clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__1159\,
            PADOUT => \N__1158\,
            PADIN => \N__1157\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_UART_TX_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1148\,
            DIN => \N__1147\,
            DOUT => \N__1146\,
            PACKAGEPIN => \o_UART_TX_wire\
        );

    \o_UART_TX_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1148\,
            PADOUT => \N__1147\,
            PADIN => \N__1146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__469\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__267\ : CascadeMux
    port map (
            O => \N__1129\,
            I => \uartTxInst.rTxState_10_0_x2_0_o2_1_0_1_cascade_\
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__1126\,
            I => \N__1123\
        );

    \I__265\ : InMux
    port map (
            O => \N__1123\,
            I => \N__1116\
        );

    \I__264\ : InMux
    port map (
            O => \N__1122\,
            I => \N__1116\
        );

    \I__263\ : InMux
    port map (
            O => \N__1121\,
            I => \N__1113\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1116\,
            I => \uartTxInst.un2_rclkcount_5\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__1113\,
            I => \uartTxInst.un2_rclkcount_5\
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__1108\,
            I => \uartTxInst.N_20_cascade_\
        );

    \I__259\ : InMux
    port map (
            O => \N__1105\,
            I => \N__1099\
        );

    \I__258\ : InMux
    port map (
            O => \N__1104\,
            I => \N__1099\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1099\,
            I => \uartTxInst.rBitIndexZ0Z_2\
        );

    \I__256\ : CascadeMux
    port map (
            O => \N__1096\,
            I => \N__1093\
        );

    \I__255\ : InMux
    port map (
            O => \N__1093\,
            I => \N__1084\
        );

    \I__254\ : InMux
    port map (
            O => \N__1092\,
            I => \N__1081\
        );

    \I__253\ : InMux
    port map (
            O => \N__1091\,
            I => \N__1074\
        );

    \I__252\ : InMux
    port map (
            O => \N__1090\,
            I => \N__1074\
        );

    \I__251\ : InMux
    port map (
            O => \N__1089\,
            I => \N__1074\
        );

    \I__250\ : InMux
    port map (
            O => \N__1088\,
            I => \N__1071\
        );

    \I__249\ : InMux
    port map (
            O => \N__1087\,
            I => \N__1068\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1084\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1081\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1074\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1071\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1068\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__1057\,
            I => \uartTxInst.rTxState_10_0_i_a2_0_1_0_cascade_\
        );

    \I__242\ : InMux
    port map (
            O => \N__1054\,
            I => \N__1048\
        );

    \I__241\ : InMux
    port map (
            O => \N__1053\,
            I => \N__1045\
        );

    \I__240\ : InMux
    port map (
            O => \N__1052\,
            I => \N__1042\
        );

    \I__239\ : InMux
    port map (
            O => \N__1051\,
            I => \N__1039\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1048\,
            I => \N__1036\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1045\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__1042\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1039\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__234\ : Odrv4
    port map (
            O => \N__1036\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__233\ : CascadeMux
    port map (
            O => \N__1027\,
            I => \N__1020\
        );

    \I__232\ : InMux
    port map (
            O => \N__1026\,
            I => \N__1014\
        );

    \I__231\ : InMux
    port map (
            O => \N__1025\,
            I => \N__1005\
        );

    \I__230\ : InMux
    port map (
            O => \N__1024\,
            I => \N__1005\
        );

    \I__229\ : InMux
    port map (
            O => \N__1023\,
            I => \N__1005\
        );

    \I__228\ : InMux
    port map (
            O => \N__1020\,
            I => \N__1005\
        );

    \I__227\ : InMux
    port map (
            O => \N__1019\,
            I => \N__1000\
        );

    \I__226\ : InMux
    port map (
            O => \N__1018\,
            I => \N__1000\
        );

    \I__225\ : InMux
    port map (
            O => \N__1017\,
            I => \N__997\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__1014\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1005\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1000\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__997\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__220\ : CascadeMux
    port map (
            O => \N__988\,
            I => \N__981\
        );

    \I__219\ : InMux
    port map (
            O => \N__987\,
            I => \N__978\
        );

    \I__218\ : InMux
    port map (
            O => \N__986\,
            I => \N__969\
        );

    \I__217\ : InMux
    port map (
            O => \N__985\,
            I => \N__969\
        );

    \I__216\ : InMux
    port map (
            O => \N__984\,
            I => \N__969\
        );

    \I__215\ : InMux
    port map (
            O => \N__981\,
            I => \N__969\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__978\,
            I => \uartTxInst.rBitIndexZ1Z_0\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__969\,
            I => \uartTxInst.rBitIndexZ1Z_0\
        );

    \I__212\ : CascadeMux
    port map (
            O => \N__964\,
            I => \N__961\
        );

    \I__211\ : InMux
    port map (
            O => \N__961\,
            I => \N__950\
        );

    \I__210\ : InMux
    port map (
            O => \N__960\,
            I => \N__941\
        );

    \I__209\ : InMux
    port map (
            O => \N__959\,
            I => \N__941\
        );

    \I__208\ : InMux
    port map (
            O => \N__958\,
            I => \N__941\
        );

    \I__207\ : InMux
    port map (
            O => \N__957\,
            I => \N__941\
        );

    \I__206\ : InMux
    port map (
            O => \N__956\,
            I => \N__936\
        );

    \I__205\ : InMux
    port map (
            O => \N__955\,
            I => \N__936\
        );

    \I__204\ : InMux
    port map (
            O => \N__954\,
            I => \N__931\
        );

    \I__203\ : InMux
    port map (
            O => \N__953\,
            I => \N__931\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__950\,
            I => \uartTxInst.rClkCountZ0Z_0\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__941\,
            I => \uartTxInst.rClkCountZ0Z_0\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__936\,
            I => \uartTxInst.rClkCountZ0Z_0\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__931\,
            I => \uartTxInst.rClkCountZ0Z_0\
        );

    \I__198\ : InMux
    port map (
            O => \N__922\,
            I => \N__919\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__919\,
            I => \uartTxInst.rBitIndex_RNO_2Z0Z_1\
        );

    \I__196\ : InMux
    port map (
            O => \N__916\,
            I => \N__911\
        );

    \I__195\ : InMux
    port map (
            O => \N__915\,
            I => \N__908\
        );

    \I__194\ : InMux
    port map (
            O => \N__914\,
            I => \N__905\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__911\,
            I => \uartTxInst.un2_rclkcount_4\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__908\,
            I => \uartTxInst.un2_rclkcount_4\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__905\,
            I => \uartTxInst.un2_rclkcount_4\
        );

    \I__190\ : CascadeMux
    port map (
            O => \N__898\,
            I => \N__886\
        );

    \I__189\ : SRMux
    port map (
            O => \N__897\,
            I => \N__881\
        );

    \I__188\ : SRMux
    port map (
            O => \N__896\,
            I => \N__878\
        );

    \I__187\ : InMux
    port map (
            O => \N__895\,
            I => \N__873\
        );

    \I__186\ : InMux
    port map (
            O => \N__894\,
            I => \N__873\
        );

    \I__185\ : InMux
    port map (
            O => \N__893\,
            I => \N__864\
        );

    \I__184\ : InMux
    port map (
            O => \N__892\,
            I => \N__864\
        );

    \I__183\ : InMux
    port map (
            O => \N__891\,
            I => \N__864\
        );

    \I__182\ : InMux
    port map (
            O => \N__890\,
            I => \N__864\
        );

    \I__181\ : InMux
    port map (
            O => \N__889\,
            I => \N__859\
        );

    \I__180\ : InMux
    port map (
            O => \N__886\,
            I => \N__859\
        );

    \I__179\ : InMux
    port map (
            O => \N__885\,
            I => \N__854\
        );

    \I__178\ : InMux
    port map (
            O => \N__884\,
            I => \N__854\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__881\,
            I => \uartTxInst.rbitindex15\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__878\,
            I => \uartTxInst.rbitindex15\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__873\,
            I => \uartTxInst.rbitindex15\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__864\,
            I => \uartTxInst.rbitindex15\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__859\,
            I => \uartTxInst.rbitindex15\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__854\,
            I => \uartTxInst.rbitindex15\
        );

    \I__171\ : CascadeMux
    port map (
            O => \N__841\,
            I => \uartTxInst.SUM_i_o2_d_1_cascade_\
        );

    \I__170\ : InMux
    port map (
            O => \N__838\,
            I => \N__835\
        );

    \I__169\ : LocalMux
    port map (
            O => \N__835\,
            I => \uartTxInst.SUM_i_o2_1_0_1\
        );

    \I__168\ : InMux
    port map (
            O => \N__832\,
            I => \N__823\
        );

    \I__167\ : InMux
    port map (
            O => \N__831\,
            I => \N__823\
        );

    \I__166\ : InMux
    port map (
            O => \N__830\,
            I => \N__823\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__823\,
            I => \uartTxInst.rBitIndexZ0Z_1\
        );

    \I__164\ : ClkMux
    port map (
            O => \N__820\,
            I => \N__802\
        );

    \I__163\ : ClkMux
    port map (
            O => \N__819\,
            I => \N__802\
        );

    \I__162\ : ClkMux
    port map (
            O => \N__818\,
            I => \N__802\
        );

    \I__161\ : ClkMux
    port map (
            O => \N__817\,
            I => \N__802\
        );

    \I__160\ : ClkMux
    port map (
            O => \N__816\,
            I => \N__802\
        );

    \I__159\ : ClkMux
    port map (
            O => \N__815\,
            I => \N__802\
        );

    \I__158\ : GlobalMux
    port map (
            O => \N__802\,
            I => \N__799\
        );

    \I__157\ : gio2CtrlBuf
    port map (
            O => \N__799\,
            I => \i_Clk_c_g\
        );

    \I__156\ : InMux
    port map (
            O => \N__796\,
            I => \N__793\
        );

    \I__155\ : LocalMux
    port map (
            O => \N__793\,
            I => \uartTxInst.N_17_mux\
        );

    \I__154\ : CascadeMux
    port map (
            O => \N__790\,
            I => \N__782\
        );

    \I__153\ : InMux
    port map (
            O => \N__789\,
            I => \N__777\
        );

    \I__152\ : InMux
    port map (
            O => \N__788\,
            I => \N__774\
        );

    \I__151\ : InMux
    port map (
            O => \N__787\,
            I => \N__767\
        );

    \I__150\ : InMux
    port map (
            O => \N__786\,
            I => \N__767\
        );

    \I__149\ : InMux
    port map (
            O => \N__785\,
            I => \N__767\
        );

    \I__148\ : InMux
    port map (
            O => \N__782\,
            I => \N__764\
        );

    \I__147\ : InMux
    port map (
            O => \N__781\,
            I => \N__759\
        );

    \I__146\ : InMux
    port map (
            O => \N__780\,
            I => \N__759\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__777\,
            I => \uartTxInst.rClkCountZ0Z_1\
        );

    \I__144\ : LocalMux
    port map (
            O => \N__774\,
            I => \uartTxInst.rClkCountZ0Z_1\
        );

    \I__143\ : LocalMux
    port map (
            O => \N__767\,
            I => \uartTxInst.rClkCountZ0Z_1\
        );

    \I__142\ : LocalMux
    port map (
            O => \N__764\,
            I => \uartTxInst.rClkCountZ0Z_1\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__759\,
            I => \uartTxInst.rClkCountZ0Z_1\
        );

    \I__140\ : CascadeMux
    port map (
            O => \N__748\,
            I => \N__743\
        );

    \I__139\ : CascadeMux
    port map (
            O => \N__747\,
            I => \N__736\
        );

    \I__138\ : InMux
    port map (
            O => \N__746\,
            I => \N__727\
        );

    \I__137\ : InMux
    port map (
            O => \N__743\,
            I => \N__727\
        );

    \I__136\ : InMux
    port map (
            O => \N__742\,
            I => \N__727\
        );

    \I__135\ : InMux
    port map (
            O => \N__741\,
            I => \N__727\
        );

    \I__134\ : InMux
    port map (
            O => \N__740\,
            I => \N__724\
        );

    \I__133\ : InMux
    port map (
            O => \N__739\,
            I => \N__719\
        );

    \I__132\ : InMux
    port map (
            O => \N__736\,
            I => \N__719\
        );

    \I__131\ : LocalMux
    port map (
            O => \N__727\,
            I => \uartTxInst.rClkCountZ0Z_2\
        );

    \I__130\ : LocalMux
    port map (
            O => \N__724\,
            I => \uartTxInst.rClkCountZ0Z_2\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__719\,
            I => \uartTxInst.rClkCountZ0Z_2\
        );

    \I__128\ : CascadeMux
    port map (
            O => \N__712\,
            I => \N__703\
        );

    \I__127\ : CascadeMux
    port map (
            O => \N__711\,
            I => \N__700\
        );

    \I__126\ : InMux
    port map (
            O => \N__710\,
            I => \N__695\
        );

    \I__125\ : InMux
    port map (
            O => \N__709\,
            I => \N__695\
        );

    \I__124\ : InMux
    port map (
            O => \N__708\,
            I => \N__688\
        );

    \I__123\ : InMux
    port map (
            O => \N__707\,
            I => \N__688\
        );

    \I__122\ : InMux
    port map (
            O => \N__706\,
            I => \N__688\
        );

    \I__121\ : InMux
    port map (
            O => \N__703\,
            I => \N__683\
        );

    \I__120\ : InMux
    port map (
            O => \N__700\,
            I => \N__683\
        );

    \I__119\ : LocalMux
    port map (
            O => \N__695\,
            I => \N__680\
        );

    \I__118\ : LocalMux
    port map (
            O => \N__688\,
            I => \uartTxInst.rClkCountZ0Z_5\
        );

    \I__117\ : LocalMux
    port map (
            O => \N__683\,
            I => \uartTxInst.rClkCountZ0Z_5\
        );

    \I__116\ : Odrv4
    port map (
            O => \N__680\,
            I => \uartTxInst.rClkCountZ0Z_5\
        );

    \I__115\ : CascadeMux
    port map (
            O => \N__673\,
            I => \uartTxInst.un2_rclkcount_5_cascade_\
        );

    \I__114\ : InMux
    port map (
            O => \N__670\,
            I => \N__667\
        );

    \I__113\ : LocalMux
    port map (
            O => \N__667\,
            I => \uartTxInst.rClkCount_RNIOIKC_0Z0Z_3\
        );

    \I__112\ : CascadeMux
    port map (
            O => \N__664\,
            I => \uartTxInst.SUM_N_3_mux_cascade_\
        );

    \I__111\ : CascadeMux
    port map (
            O => \N__661\,
            I => \N__657\
        );

    \I__110\ : InMux
    port map (
            O => \N__660\,
            I => \N__653\
        );

    \I__109\ : InMux
    port map (
            O => \N__657\,
            I => \N__648\
        );

    \I__108\ : InMux
    port map (
            O => \N__656\,
            I => \N__648\
        );

    \I__107\ : LocalMux
    port map (
            O => \N__653\,
            I => \uartTxInst.un5_rclkcount_c4\
        );

    \I__106\ : LocalMux
    port map (
            O => \N__648\,
            I => \uartTxInst.un5_rclkcount_c4\
        );

    \I__105\ : CascadeMux
    port map (
            O => \N__643\,
            I => \N__638\
        );

    \I__104\ : CascadeMux
    port map (
            O => \N__642\,
            I => \N__632\
        );

    \I__103\ : InMux
    port map (
            O => \N__641\,
            I => \N__627\
        );

    \I__102\ : InMux
    port map (
            O => \N__638\,
            I => \N__622\
        );

    \I__101\ : InMux
    port map (
            O => \N__637\,
            I => \N__622\
        );

    \I__100\ : InMux
    port map (
            O => \N__636\,
            I => \N__617\
        );

    \I__99\ : InMux
    port map (
            O => \N__635\,
            I => \N__617\
        );

    \I__98\ : InMux
    port map (
            O => \N__632\,
            I => \N__610\
        );

    \I__97\ : InMux
    port map (
            O => \N__631\,
            I => \N__610\
        );

    \I__96\ : InMux
    port map (
            O => \N__630\,
            I => \N__610\
        );

    \I__95\ : LocalMux
    port map (
            O => \N__627\,
            I => \uartTxInst.rClkCountZ0Z_4\
        );

    \I__94\ : LocalMux
    port map (
            O => \N__622\,
            I => \uartTxInst.rClkCountZ0Z_4\
        );

    \I__93\ : LocalMux
    port map (
            O => \N__617\,
            I => \uartTxInst.rClkCountZ0Z_4\
        );

    \I__92\ : LocalMux
    port map (
            O => \N__610\,
            I => \uartTxInst.rClkCountZ0Z_4\
        );

    \I__91\ : InMux
    port map (
            O => \N__601\,
            I => \N__592\
        );

    \I__90\ : InMux
    port map (
            O => \N__600\,
            I => \N__592\
        );

    \I__89\ : InMux
    port map (
            O => \N__599\,
            I => \N__589\
        );

    \I__88\ : InMux
    port map (
            O => \N__598\,
            I => \N__584\
        );

    \I__87\ : InMux
    port map (
            O => \N__597\,
            I => \N__584\
        );

    \I__86\ : LocalMux
    port map (
            O => \N__592\,
            I => \uartTxInst.rClkCountZ0Z_3\
        );

    \I__85\ : LocalMux
    port map (
            O => \N__589\,
            I => \uartTxInst.rClkCountZ0Z_3\
        );

    \I__84\ : LocalMux
    port map (
            O => \N__584\,
            I => \uartTxInst.rClkCountZ0Z_3\
        );

    \I__83\ : CascadeMux
    port map (
            O => \N__577\,
            I => \N__572\
        );

    \I__82\ : InMux
    port map (
            O => \N__576\,
            I => \N__569\
        );

    \I__81\ : CascadeMux
    port map (
            O => \N__575\,
            I => \N__566\
        );

    \I__80\ : InMux
    port map (
            O => \N__572\,
            I => \N__561\
        );

    \I__79\ : LocalMux
    port map (
            O => \N__569\,
            I => \N__558\
        );

    \I__78\ : InMux
    port map (
            O => \N__566\,
            I => \N__555\
        );

    \I__77\ : InMux
    port map (
            O => \N__565\,
            I => \N__550\
        );

    \I__76\ : InMux
    port map (
            O => \N__564\,
            I => \N__550\
        );

    \I__75\ : LocalMux
    port map (
            O => \N__561\,
            I => \uartTxInst.rClkCountZ0Z_7\
        );

    \I__74\ : Odrv4
    port map (
            O => \N__558\,
            I => \uartTxInst.rClkCountZ0Z_7\
        );

    \I__73\ : LocalMux
    port map (
            O => \N__555\,
            I => \uartTxInst.rClkCountZ0Z_7\
        );

    \I__72\ : LocalMux
    port map (
            O => \N__550\,
            I => \uartTxInst.rClkCountZ0Z_7\
        );

    \I__71\ : CascadeMux
    port map (
            O => \N__541\,
            I => \N__533\
        );

    \I__70\ : InMux
    port map (
            O => \N__540\,
            I => \N__528\
        );

    \I__69\ : InMux
    port map (
            O => \N__539\,
            I => \N__528\
        );

    \I__68\ : InMux
    port map (
            O => \N__538\,
            I => \N__523\
        );

    \I__67\ : InMux
    port map (
            O => \N__537\,
            I => \N__523\
        );

    \I__66\ : InMux
    port map (
            O => \N__536\,
            I => \N__520\
        );

    \I__65\ : InMux
    port map (
            O => \N__533\,
            I => \N__517\
        );

    \I__64\ : LocalMux
    port map (
            O => \N__528\,
            I => \uartTxInst.rClkCountZ0Z_6\
        );

    \I__63\ : LocalMux
    port map (
            O => \N__523\,
            I => \uartTxInst.rClkCountZ0Z_6\
        );

    \I__62\ : LocalMux
    port map (
            O => \N__520\,
            I => \uartTxInst.rClkCountZ0Z_6\
        );

    \I__61\ : LocalMux
    port map (
            O => \N__517\,
            I => \uartTxInst.rClkCountZ0Z_6\
        );

    \I__60\ : CascadeMux
    port map (
            O => \N__508\,
            I => \uartTxInst.un2_rclkcount_4_cascade_\
        );

    \I__59\ : CascadeMux
    port map (
            O => \N__505\,
            I => \uartTxInst.un5_rclkcount_ac0_11_cascade_\
        );

    \I__58\ : CascadeMux
    port map (
            O => \N__502\,
            I => \uartTxInst.un5_rclkcount_c4_cascade_\
        );

    \I__57\ : CascadeMux
    port map (
            O => \N__499\,
            I => \uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_\
        );

    \I__56\ : CascadeMux
    port map (
            O => \N__496\,
            I => \uartTxInst.N_8_i_cascade_\
        );

    \I__55\ : InMux
    port map (
            O => \N__493\,
            I => \N__490\
        );

    \I__54\ : LocalMux
    port map (
            O => \N__490\,
            I => \uartTxInst.m11_i_a3_3\
        );

    \I__53\ : InMux
    port map (
            O => \N__487\,
            I => \N__484\
        );

    \I__52\ : LocalMux
    port map (
            O => \N__484\,
            I => \uartTxInst.m11_i_a3_4\
        );

    \I__51\ : InMux
    port map (
            O => \N__481\,
            I => \N__478\
        );

    \I__50\ : LocalMux
    port map (
            O => \N__478\,
            I => \uartTxInst.m15_e_5\
        );

    \I__49\ : InMux
    port map (
            O => \N__475\,
            I => \N__472\
        );

    \I__48\ : LocalMux
    port map (
            O => \N__472\,
            I => \uartTxInst.m15_e_4\
        );

    \I__47\ : IoInMux
    port map (
            O => \N__469\,
            I => \N__466\
        );

    \I__46\ : LocalMux
    port map (
            O => \N__466\,
            I => \N__463\
        );

    \I__45\ : IoSpan4Mux
    port map (
            O => \N__463\,
            I => \N__460\
        );

    \I__44\ : Span4Mux_s3_h
    port map (
            O => \N__460\,
            I => \N__456\
        );

    \I__43\ : CascadeMux
    port map (
            O => \N__459\,
            I => \N__453\
        );

    \I__42\ : Span4Mux_h
    port map (
            O => \N__456\,
            I => \N__450\
        );

    \I__41\ : InMux
    port map (
            O => \N__453\,
            I => \N__447\
        );

    \I__40\ : Odrv4
    port map (
            O => \N__450\,
            I => \o_UART_TX_c\
        );

    \I__39\ : LocalMux
    port map (
            O => \N__447\,
            I => \o_UART_TX_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNO_0_3_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101010101"
        )
    port map (
            in0 => \N__601\,
            in1 => \N__787\,
            in2 => \N__748\,
            in3 => \N__959\,
            lcout => OPEN,
            ltout => \uartTxInst.N_8_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_3_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__889\,
            in1 => \N__487\,
            in2 => \N__496\,
            in3 => \N__493\,
            lcout => \uartTxInst.rClkCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNO_1_3_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__576\,
            in1 => \_gnd_net_\,
            in2 => \N__712\,
            in3 => \N__957\,
            lcout => \uartTxInst.m11_i_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_2_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__960\,
            in1 => \N__746\,
            in2 => \N__898\,
            in3 => \N__789\,
            lcout => \uartTxInst.rClkCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.oSerial_RNO_1_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__741\,
            in1 => \N__785\,
            in2 => \N__711\,
            in3 => \N__958\,
            lcout => \uartTxInst.m15_e_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNO_2_3_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__742\,
            in1 => \N__538\,
            in2 => \N__643\,
            in3 => \N__786\,
            lcout => \uartTxInst.m11_i_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.oSerial_RNO_2_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__537\,
            in1 => \N__637\,
            in2 => \N__577\,
            in3 => \N__600\,
            lcout => \uartTxInst.m15_e_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.oSerial_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__481\,
            in1 => \N__475\,
            in2 => \N__459\,
            in3 => \N__796\,
            lcout => \o_UART_TX_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__816\,
            ce => 'H',
            sr => \N__896\
        );

    \uartTxInst.rTxState_RNINSDP_1_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1088\,
            in2 => \_gnd_net_\,
            in3 => \N__1017\,
            lcout => \uartTxInst.rbitindex15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_0_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001001"
        )
    port map (
            in0 => \N__1026\,
            in1 => \N__987\,
            in2 => \N__1096\,
            in3 => \N__1052\,
            lcout => \uartTxInst.rBitIndexZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__818\,
            ce => 'H',
            sr => \N__897\
        );

    \uartTxInst.rClkCount_RNO_0_7_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__706\,
            in1 => \N__539\,
            in2 => \N__642\,
            in3 => \N__656\,
            lcout => OPEN,
            ltout => \uartTxInst.un5_rclkcount_ac0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_7_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__565\,
            in1 => \N__892\,
            in2 => \N__505\,
            in3 => \N__1053\,
            lcout => \uartTxInst.rClkCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNIOIKC_0_3_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__630\,
            in1 => \N__597\,
            in2 => \N__541\,
            in3 => \N__564\,
            lcout => \uartTxInst.rClkCount_RNIOIKC_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_5_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__641\,
            in1 => \N__891\,
            in2 => \N__661\,
            in3 => \N__708\,
            lcout => \uartTxInst.rClkCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNIA4KC_3_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__955\,
            in1 => \N__598\,
            in2 => \N__790\,
            in3 => \N__740\,
            lcout => \uartTxInst.un5_rclkcount_c4\,
            ltout => \uartTxInst.un5_rclkcount_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNO_0_6_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__540\,
            in1 => \N__631\,
            in2 => \N__502\,
            in3 => \N__707\,
            lcout => OPEN,
            ltout => \uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_6_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__893\,
            in1 => \_gnd_net_\,
            in2 => \N__499\,
            in3 => \N__1054\,
            lcout => \uartTxInst.rClkCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__788\,
            in1 => \N__956\,
            in2 => \_gnd_net_\,
            in3 => \N__890\,
            lcout => \uartTxInst.rClkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__954\,
            in1 => \N__884\,
            in2 => \N__1126\,
            in3 => \N__916\,
            lcout => \uartTxInst.rClkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.oSerial_RNO_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1087\,
            in2 => \_gnd_net_\,
            in3 => \N__1018\,
            lcout => \uartTxInst.N_17_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNO_2_1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__710\,
            in1 => \N__739\,
            in2 => \_gnd_net_\,
            in3 => \N__781\,
            lcout => \uartTxInst.rBitIndex_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNIC6KC_2_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__780\,
            in1 => \N__953\,
            in2 => \N__747\,
            in3 => \N__709\,
            lcout => \uartTxInst.un2_rclkcount_5\,
            ltout => \uartTxInst.un2_rclkcount_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNI4P8P_3_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__673\,
            in3 => \N__670\,
            lcout => \uartTxInst.SUM_N_3_mux\,
            ltout => \uartTxInst.SUM_N_3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_4_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__885\,
            in1 => \N__636\,
            in2 => \N__664\,
            in3 => \N__660\,
            lcout => \uartTxInst.rClkCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNIOIKC_3_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__635\,
            in1 => \N__599\,
            in2 => \N__575\,
            in3 => \N__536\,
            lcout => \uartTxInst.un2_rclkcount_4\,
            ltout => \uartTxInst.un2_rclkcount_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxState_1_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__1092\,
            in1 => \N__1019\,
            in2 => \N__508\,
            in3 => \N__1122\,
            lcout => \uartTxInst.rTxStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNO_0_1_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010101"
        )
    port map (
            in0 => \N__831\,
            in1 => \N__1089\,
            in2 => \N__1027\,
            in3 => \N__984\,
            lcout => \uartTxInst.SUM_i_o2_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNO_1_2_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1023\,
            in2 => \N__988\,
            in3 => \N__830\,
            lcout => OPEN,
            ltout => \uartTxInst.rTxState_10_0_x2_0_o2_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNO_0_2_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111100"
        )
    port map (
            in0 => \N__914\,
            in1 => \N__1090\,
            in2 => \N__1129\,
            in3 => \N__1121\,
            lcout => OPEN,
            ltout => \uartTxInst.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_2_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100101"
        )
    port map (
            in0 => \N__1105\,
            in1 => \_gnd_net_\,
            in2 => \N__1108\,
            in3 => \N__894\,
            lcout => \uartTxInst.rBitIndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxState_RNO_0_0_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__832\,
            in1 => \N__1104\,
            in2 => \_gnd_net_\,
            in3 => \N__1091\,
            lcout => OPEN,
            ltout => \uartTxInst.rTxState_10_0_i_a2_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxState_0_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000011001100"
        )
    port map (
            in0 => \N__986\,
            in1 => \N__1025\,
            in2 => \N__1057\,
            in3 => \N__1051\,
            lcout => \uartTxInst.rTxStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNO_1_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__1024\,
            in1 => \N__985\,
            in2 => \N__964\,
            in3 => \N__922\,
            lcout => OPEN,
            ltout => \uartTxInst.SUM_i_o2_d_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_1_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000110001"
        )
    port map (
            in0 => \N__915\,
            in1 => \N__895\,
            in2 => \N__841\,
            in3 => \N__838\,
            lcout => \uartTxInst.rBitIndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__820\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
