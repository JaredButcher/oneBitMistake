// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 28 2019 14:20:42

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "core" view "INTERFACE"

module core (
    o_UART_TX,
    i_UART_RX,
    i_Clk);

    output o_UART_TX;
    input i_UART_RX;
    input i_Clk;

    wire N__3127;
    wire N__3126;
    wire N__3125;
    wire N__3116;
    wire N__3115;
    wire N__3114;
    wire N__3107;
    wire N__3106;
    wire N__3105;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3081;
    wire N__3078;
    wire N__3077;
    wire N__3076;
    wire N__3075;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3052;
    wire N__3051;
    wire N__3050;
    wire N__3049;
    wire N__3048;
    wire N__3047;
    wire N__3046;
    wire N__3045;
    wire N__3044;
    wire N__3043;
    wire N__3042;
    wire N__3041;
    wire N__3040;
    wire N__3037;
    wire N__3028;
    wire N__3025;
    wire N__3020;
    wire N__3015;
    wire N__3008;
    wire N__3003;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2982;
    wire N__2981;
    wire N__2980;
    wire N__2979;
    wire N__2978;
    wire N__2973;
    wire N__2972;
    wire N__2969;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2942;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2926;
    wire N__2925;
    wire N__2924;
    wire N__2923;
    wire N__2922;
    wire N__2919;
    wire N__2918;
    wire N__2917;
    wire N__2916;
    wire N__2911;
    wire N__2910;
    wire N__2909;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2901;
    wire N__2898;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2882;
    wire N__2873;
    wire N__2860;
    wire N__2857;
    wire N__2854;
    wire N__2851;
    wire N__2850;
    wire N__2849;
    wire N__2848;
    wire N__2847;
    wire N__2846;
    wire N__2845;
    wire N__2842;
    wire N__2835;
    wire N__2828;
    wire N__2821;
    wire N__2820;
    wire N__2819;
    wire N__2818;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2804;
    wire N__2797;
    wire N__2796;
    wire N__2795;
    wire N__2794;
    wire N__2793;
    wire N__2792;
    wire N__2791;
    wire N__2790;
    wire N__2789;
    wire N__2788;
    wire N__2787;
    wire N__2786;
    wire N__2785;
    wire N__2784;
    wire N__2783;
    wire N__2782;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2735;
    wire N__2732;
    wire N__2729;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2710;
    wire N__2709;
    wire N__2708;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire N__2696;
    wire N__2689;
    wire N__2686;
    wire N__2685;
    wire N__2684;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2674;
    wire N__2671;
    wire N__2662;
    wire N__2661;
    wire N__2660;
    wire N__2657;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2647;
    wire N__2642;
    wire N__2635;
    wire N__2634;
    wire N__2633;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2611;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2580;
    wire N__2577;
    wire N__2574;
    wire N__2569;
    wire N__2566;
    wire N__2563;
    wire N__2560;
    wire N__2557;
    wire N__2554;
    wire N__2551;
    wire N__2548;
    wire N__2547;
    wire N__2546;
    wire N__2545;
    wire N__2544;
    wire N__2541;
    wire N__2538;
    wire N__2531;
    wire N__2528;
    wire N__2521;
    wire N__2520;
    wire N__2519;
    wire N__2518;
    wire N__2517;
    wire N__2514;
    wire N__2509;
    wire N__2504;
    wire N__2497;
    wire N__2494;
    wire N__2493;
    wire N__2492;
    wire N__2491;
    wire N__2488;
    wire N__2481;
    wire N__2476;
    wire N__2473;
    wire N__2472;
    wire N__2467;
    wire N__2464;
    wire N__2463;
    wire N__2460;
    wire N__2459;
    wire N__2452;
    wire N__2449;
    wire N__2446;
    wire N__2443;
    wire N__2442;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2430;
    wire N__2425;
    wire N__2422;
    wire N__2419;
    wire N__2416;
    wire N__2413;
    wire N__2412;
    wire N__2409;
    wire N__2406;
    wire N__2401;
    wire N__2398;
    wire N__2397;
    wire N__2394;
    wire N__2391;
    wire N__2386;
    wire N__2383;
    wire N__2382;
    wire N__2379;
    wire N__2376;
    wire N__2371;
    wire N__2368;
    wire N__2365;
    wire N__2362;
    wire N__2359;
    wire N__2356;
    wire N__2353;
    wire N__2350;
    wire N__2347;
    wire N__2344;
    wire N__2341;
    wire N__2338;
    wire N__2335;
    wire N__2332;
    wire N__2329;
    wire N__2326;
    wire N__2323;
    wire N__2320;
    wire N__2317;
    wire N__2314;
    wire N__2311;
    wire N__2308;
    wire N__2305;
    wire N__2304;
    wire N__2301;
    wire N__2300;
    wire N__2299;
    wire N__2298;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2288;
    wire N__2285;
    wire N__2282;
    wire N__2279;
    wire N__2276;
    wire N__2263;
    wire N__2260;
    wire N__2257;
    wire N__2254;
    wire N__2253;
    wire N__2252;
    wire N__2249;
    wire N__2246;
    wire N__2243;
    wire N__2236;
    wire N__2233;
    wire N__2230;
    wire N__2227;
    wire N__2224;
    wire N__2221;
    wire N__2220;
    wire N__2217;
    wire N__2214;
    wire N__2209;
    wire N__2206;
    wire N__2205;
    wire N__2202;
    wire N__2199;
    wire N__2194;
    wire N__2191;
    wire N__2188;
    wire N__2185;
    wire N__2184;
    wire N__2181;
    wire N__2178;
    wire N__2173;
    wire N__2170;
    wire N__2169;
    wire N__2166;
    wire N__2163;
    wire N__2158;
    wire N__2155;
    wire N__2152;
    wire N__2149;
    wire N__2146;
    wire N__2145;
    wire N__2142;
    wire N__2139;
    wire N__2134;
    wire N__2131;
    wire N__2130;
    wire N__2127;
    wire N__2124;
    wire N__2119;
    wire N__2116;
    wire N__2113;
    wire N__2110;
    wire N__2107;
    wire N__2104;
    wire N__2103;
    wire N__2100;
    wire N__2099;
    wire N__2096;
    wire N__2091;
    wire N__2086;
    wire N__2083;
    wire N__2082;
    wire N__2081;
    wire N__2080;
    wire N__2077;
    wire N__2070;
    wire N__2065;
    wire N__2062;
    wire N__2059;
    wire N__2056;
    wire N__2053;
    wire N__2050;
    wire N__2047;
    wire N__2044;
    wire N__2041;
    wire N__2038;
    wire N__2035;
    wire N__2032;
    wire N__2031;
    wire N__2030;
    wire N__2027;
    wire N__2024;
    wire N__2021;
    wire N__2020;
    wire N__2019;
    wire N__2018;
    wire N__2011;
    wire N__2010;
    wire N__2009;
    wire N__2006;
    wire N__2003;
    wire N__2000;
    wire N__1997;
    wire N__1994;
    wire N__1991;
    wire N__1984;
    wire N__1979;
    wire N__1976;
    wire N__1973;
    wire N__1970;
    wire N__1967;
    wire N__1960;
    wire N__1957;
    wire N__1954;
    wire N__1951;
    wire N__1950;
    wire N__1949;
    wire N__1948;
    wire N__1943;
    wire N__1940;
    wire N__1937;
    wire N__1930;
    wire N__1929;
    wire N__1926;
    wire N__1923;
    wire N__1920;
    wire N__1915;
    wire N__1914;
    wire N__1911;
    wire N__1908;
    wire N__1903;
    wire N__1902;
    wire N__1901;
    wire N__1900;
    wire N__1899;
    wire N__1896;
    wire N__1893;
    wire N__1890;
    wire N__1885;
    wire N__1882;
    wire N__1873;
    wire N__1872;
    wire N__1869;
    wire N__1866;
    wire N__1861;
    wire N__1858;
    wire N__1855;
    wire N__1854;
    wire N__1851;
    wire N__1848;
    wire N__1843;
    wire N__1842;
    wire N__1841;
    wire N__1838;
    wire N__1835;
    wire N__1832;
    wire N__1825;
    wire N__1822;
    wire N__1821;
    wire N__1820;
    wire N__1819;
    wire N__1818;
    wire N__1817;
    wire N__1816;
    wire N__1815;
    wire N__1812;
    wire N__1809;
    wire N__1806;
    wire N__1797;
    wire N__1794;
    wire N__1783;
    wire N__1780;
    wire N__1777;
    wire N__1774;
    wire N__1773;
    wire N__1768;
    wire N__1765;
    wire N__1762;
    wire N__1759;
    wire N__1756;
    wire N__1755;
    wire N__1754;
    wire N__1751;
    wire N__1750;
    wire N__1749;
    wire N__1746;
    wire N__1743;
    wire N__1742;
    wire N__1741;
    wire N__1740;
    wire N__1739;
    wire N__1734;
    wire N__1731;
    wire N__1722;
    wire N__1717;
    wire N__1708;
    wire N__1705;
    wire N__1702;
    wire N__1699;
    wire N__1696;
    wire N__1693;
    wire N__1690;
    wire N__1689;
    wire N__1686;
    wire N__1683;
    wire N__1678;
    wire N__1677;
    wire N__1676;
    wire N__1673;
    wire N__1672;
    wire N__1671;
    wire N__1670;
    wire N__1669;
    wire N__1668;
    wire N__1667;
    wire N__1666;
    wire N__1665;
    wire N__1662;
    wire N__1661;
    wire N__1660;
    wire N__1657;
    wire N__1656;
    wire N__1653;
    wire N__1650;
    wire N__1639;
    wire N__1632;
    wire N__1627;
    wire N__1622;
    wire N__1609;
    wire N__1608;
    wire N__1607;
    wire N__1606;
    wire N__1605;
    wire N__1602;
    wire N__1593;
    wire N__1590;
    wire N__1585;
    wire N__1582;
    wire N__1579;
    wire N__1578;
    wire N__1577;
    wire N__1574;
    wire N__1571;
    wire N__1568;
    wire N__1561;
    wire N__1560;
    wire N__1557;
    wire N__1556;
    wire N__1555;
    wire N__1552;
    wire N__1547;
    wire N__1544;
    wire N__1537;
    wire N__1536;
    wire N__1535;
    wire N__1532;
    wire N__1525;
    wire N__1522;
    wire N__1521;
    wire N__1520;
    wire N__1519;
    wire N__1518;
    wire N__1517;
    wire N__1516;
    wire N__1515;
    wire N__1514;
    wire N__1513;
    wire N__1508;
    wire N__1505;
    wire N__1500;
    wire N__1497;
    wire N__1494;
    wire N__1487;
    wire N__1484;
    wire N__1471;
    wire N__1468;
    wire N__1467;
    wire N__1466;
    wire N__1465;
    wire N__1464;
    wire N__1461;
    wire N__1458;
    wire N__1451;
    wire N__1448;
    wire N__1441;
    wire N__1438;
    wire N__1435;
    wire N__1432;
    wire N__1429;
    wire N__1426;
    wire N__1423;
    wire N__1420;
    wire N__1419;
    wire N__1416;
    wire N__1413;
    wire N__1410;
    wire N__1407;
    wire N__1402;
    wire N__1399;
    wire N__1398;
    wire N__1397;
    wire N__1396;
    wire N__1395;
    wire N__1388;
    wire N__1383;
    wire N__1378;
    wire N__1375;
    wire N__1374;
    wire N__1371;
    wire N__1368;
    wire N__1363;
    wire N__1362;
    wire N__1361;
    wire N__1356;
    wire N__1353;
    wire N__1348;
    wire N__1347;
    wire N__1346;
    wire N__1343;
    wire N__1340;
    wire N__1339;
    wire N__1338;
    wire N__1331;
    wire N__1326;
    wire N__1321;
    wire N__1320;
    wire N__1319;
    wire N__1318;
    wire N__1317;
    wire N__1316;
    wire N__1315;
    wire N__1306;
    wire N__1299;
    wire N__1294;
    wire N__1291;
    wire N__1288;
    wire N__1285;
    wire N__1282;
    wire N__1279;
    wire VCCG0;
    wire GNDG0;
    wire \uartTxInst.un5_rclkcount_c4_cascade_ ;
    wire \uartTxInst.un5_rclkcount_ac0_11_cascade_ ;
    wire \uartTxInst.un5_rclkcount_c3_cascade_ ;
    wire \uartTxInst.rbitindex15_cascade_ ;
    wire \uartTxInst.rClkCountZ0Z_1 ;
    wire \uartTxInst.un2_rclkcount_5_0_cascade_ ;
    wire \uartTxInst.rClkCountZ0Z_7 ;
    wire \uartTxInst.rClkCountZ0Z_3 ;
    wire \uartTxInst.rClkCountZ0Z_2 ;
    wire \uartTxInst.rClkCountZ0Z_0 ;
    wire \uartTxInst.un2_rclkcount_4_cascade_ ;
    wire \uartTxInst.un2_rclkcount_5_0 ;
    wire \uartTxInst.g2_0_cascade_ ;
    wire \uartTxInst.rBitIndex_RNO_0Z0Z_1_cascade_ ;
    wire \uartTxInst.rTxByte_0_sqmuxa ;
    wire \uartTxInst.rTxState_10_0_i_a2_1_2_0_cascade_ ;
    wire o_UART_TX_c;
    wire \uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_ ;
    wire \uartTxInst.rClkCountZ0Z_6 ;
    wire \uartTxInst.rClkCountZ0Z_5 ;
    wire \uartTxInst.un5_rclkcount_c4 ;
    wire \uartTxInst.SUM_N_3_mux ;
    wire \uartTxInst.rClkCountZ0Z_4 ;
    wire \uartTxInst.N_31 ;
    wire \uartTxInst.rTxStateZ0Z_1 ;
    wire \uartTxInst.un2_rclkcount_4 ;
    wire \uartTxInst.N_31_cascade_ ;
    wire \uartTxInst.rTxState_10_0_x2_0_o2_1_1_1 ;
    wire \uartTxInst.rTxState_10_0_x2_0_o2_1_1_1_cascade_ ;
    wire \uartTxInst.rTxState_10_0_x2_0_o2_d_0_1 ;
    wire \uartTxInst.rbitindex15 ;
    wire rTxDVZ0;
    wire \uartRxInst.rDataCounter_RNO_0Z0Z_1_cascade_ ;
    wire \uartTxInst.rBitIndexZ0Z_1 ;
    wire \uartTxInst.rTxByte_0_4 ;
    wire \uartTxInst.rTxByte_0_6 ;
    wire \uartTxInst.rBitIndexZ1Z_0 ;
    wire \uartTxInst.rTxByte_0_7 ;
    wire \uartTxInst.oSerial_3_6_i_m2_ns_1_cascade_ ;
    wire \uartTxInst.rTxByte_0_5 ;
    wire \uartTxInst.rBitIndexZ0Z_2 ;
    wire \uartTxInst.N_35_cascade_ ;
    wire \uartTxInst.rTxStateZ0Z_0 ;
    wire \uartTxInst.N_48 ;
    wire \uartRxInst.rDataCounterZ0Z_2 ;
    wire \uartRxInst.rstateZ0_cascade_ ;
    wire \uartRxInst.rDataCounterZ0Z_1 ;
    wire \uartRxInst.rDataCounterZ0Z_0 ;
    wire \uartRxInst.CO1_0 ;
    wire bfn_8_13_0_;
    wire \uartRxInst.rCycleCounter_cry_0 ;
    wire \uartRxInst.rCycleCounter_cry_1 ;
    wire \uartRxInst.rCycleCounter_cry_2 ;
    wire \uartRxInst.rCycleCounter_cry_3_THRU_CO ;
    wire \uartRxInst.rCycleCounter_cry_3 ;
    wire \uartRxInst.rCycleCounter_s_5 ;
    wire \uartRxInst.rCycleCounter_cry_4 ;
    wire CONSTANT_ONE_NET;
    wire \uartRxInst.rCycleCounter_s_6 ;
    wire \uartRxInst.rCycleCounter_cry_5 ;
    wire \uartRxInst.rCycleCounter_cry_6 ;
    wire rRamAddressZ0Z_0;
    wire pEcho_rRamAddress_2_0;
    wire bfn_9_9_0_;
    wire rRamAddressZ0Z_1;
    wire pEcho_rRamAddress_2_1;
    wire pEcho_rRamAddress_2_cry_0;
    wire rRamAddressZ0Z_2;
    wire pEcho_rRamAddress_2_2;
    wire pEcho_rRamAddress_2_cry_1;
    wire pEcho_rRamAddress_2_cry_2;
    wire rRamAddressZ0Z_4;
    wire pEcho_rRamAddress_2_4;
    wire pEcho_rRamAddress_2_cry_3;
    wire pEcho_rRamAddress_2_cry_4;
    wire pEcho_rRamAddress_2_5;
    wire pEcho_rRamAddress_2_5_cascade_;
    wire rRamAddressZ0Z_5;
    wire pEcho_rRamAddress_2_3;
    wire rRamAddressZ0Z_3;
    wire rRamReadData_0;
    wire rTxByteZ0Z_4;
    wire rRamReadData_1;
    wire rTxByteZ0Z_5;
    wire rRamReadData_2;
    wire rTxByteZ0Z_6;
    wire rRamReadData_3;
    wire rTxByteZ0Z_7;
    wire rRxReady;
    wire G_11_i_a3_0_6;
    wire G_11_i_a3_0_4_cascade_;
    wire uartRxInst_un1_rData_0_sqmuxa_0;
    wire N_5;
    wire \uartRxInst.un1_rCycleCounter_2_sqmuxa_0 ;
    wire \uartRxInst.rCycleCounterZ0Z_5 ;
    wire \uartRxInst.rCycleCounterZ0Z_4 ;
    wire \uartRxInst.un12_rstate_3_cascade_ ;
    wire \uartRxInst.N_83_0_i ;
    wire \uartRxInst.N_83_0_i_cascade_ ;
    wire \uartRxInst.rState_0_sqmuxa_1_1 ;
    wire \uartRxInst.rDataCounter_0_sqmuxa ;
    wire \uartRxInst.rCycleCounter_cry_0_THRU_CO ;
    wire \uartRxInst.rstateZ0 ;
    wire \uartRxInst.rCycleCounter_s_2 ;
    wire \uartRxInst.un12_rstate_4 ;
    wire \uartRxInst.rCycleCounterZ0Z_1 ;
    wire uartRxInst_rState_0;
    wire \uartRxInst.g0_0_5_cascade_ ;
    wire \uartRxInst.g0_0_4 ;
    wire i_UART_RX_c;
    wire uartRxInst_rState_1;
    wire \uartRxInst.N_83_0_i_0_cascade_ ;
    wire \uartRxInst.rCycleCounter_s_3 ;
    wire \uartRxInst.N_83_0_i_0 ;
    wire \uartRxInst.rCycleCounterZ0Z_0 ;
    wire i_Clk_c_g;
    wire \uartRxInst.rCycleCountere_0_i ;
    wire \uartRxInst.rCycleCounterZ0Z_2 ;
    wire \uartRxInst.rCycleCounterZ0Z_7 ;
    wire \uartRxInst.rCycleCounterZ0Z_3 ;
    wire \uartRxInst.rCycleCounterZ0Z_6 ;
    wire G_11_i_a3_0_5;
    wire CONSTANT_ZERO_NET;
    wire _gnd_net_;

    defparam \ramInst.rramvalues_rramvalues_0_0_physical .INIT_0=256'b0000000000000000000000000000101100000000000011110000000000000101000000000000101000000000000000000000000000001011000000000000111100000000000000000000000000001011000000000000111100000000000001010000000000001010000000000000000000000000000010110000000000001111;
    defparam \ramInst.rramvalues_rramvalues_0_0_physical .WRITE_MODE=0;
    defparam \ramInst.rramvalues_rramvalues_0_0_physical .READ_MODE=0;
    defparam \ramInst.rramvalues_rramvalues_0_0_physical .INIT_3=256'b0000000000000000000000000000101100000000000011110000000000000101000000000000101000000000000000000000000000001011000000000000111100000000000000000000000000001011000000000000111100000000000001010000000000001010000000000000000000000000000010110000000000001111;
    defparam \ramInst.rramvalues_rramvalues_0_0_physical .INIT_2=256'b0000000000000000000000000000101100000000000011110000000000000101000000000000101000000000000000000000000000001011000000000000111100000000000000000000000000001011000000000000111100000000000001010000000000001010000000000000000000000000000010110000000000001111;
    defparam \ramInst.rramvalues_rramvalues_0_0_physical .INIT_1=256'b0000000000000000000000000000101100000000000011110000000000000101000000000000101000000000000000000000000000001011000000000000111100000000000000000000000000001011000000000000111100000000000001010000000000001010000000000000000000000000000010110000000000001111;
    SB_RAM40_4K \ramInst.rramvalues_rramvalues_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,rRamReadData_3,rRamReadData_2,rRamReadData_1,rRamReadData_0}),
            .RADDR({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,N__2113,N__2134,N__2401,N__2173,N__2209,N__2236}),
            .WADDR({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,N__2416,N__2152,N__2386,N__2191,N__2227,N__2260}),
            .MASK({dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37}),
            .WDATA({dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53}),
            .RCLKE(),
            .RCLK(N__2789),
            .RE(N__2009),
            .WCLKE(N__2605),
            .WCLK(N__2790),
            .WE(N__2010));
    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3125),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__3127),
            .DIN(N__3126),
            .DOUT(N__3125),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__3127),
            .PADOUT(N__3126),
            .PADIN(N__3125),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_UART_TX_obuf_iopad (
            .OE(N__3116),
            .DIN(N__3115),
            .DOUT(N__3114),
            .PACKAGEPIN(o_UART_TX));
    defparam o_UART_TX_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_UART_TX_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_UART_TX_obuf_preio (
            .PADOEN(N__3116),
            .PADOUT(N__3115),
            .PADIN(N__3114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1426),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_UART_RX_ibuf_iopad (
            .OE(N__3107),
            .DIN(N__3106),
            .DOUT(N__3105),
            .PACKAGEPIN(i_UART_RX));
    defparam i_UART_RX_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_UART_RX_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_UART_RX_ibuf_preio (
            .PADOEN(N__3107),
            .PADOUT(N__3106),
            .PADIN(N__3105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_UART_RX_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__706 (
            .O(N__3088),
            .I(N__3085));
    LocalMux I__705 (
            .O(N__3085),
            .I(\uartRxInst.un12_rstate_4 ));
    CascadeMux I__704 (
            .O(N__3082),
            .I(N__3078));
    InMux I__703 (
            .O(N__3081),
            .I(N__3070));
    InMux I__702 (
            .O(N__3078),
            .I(N__3070));
    InMux I__701 (
            .O(N__3077),
            .I(N__3067));
    InMux I__700 (
            .O(N__3076),
            .I(N__3064));
    InMux I__699 (
            .O(N__3075),
            .I(N__3061));
    LocalMux I__698 (
            .O(N__3070),
            .I(\uartRxInst.rCycleCounterZ0Z_1 ));
    LocalMux I__697 (
            .O(N__3067),
            .I(\uartRxInst.rCycleCounterZ0Z_1 ));
    LocalMux I__696 (
            .O(N__3064),
            .I(\uartRxInst.rCycleCounterZ0Z_1 ));
    LocalMux I__695 (
            .O(N__3061),
            .I(\uartRxInst.rCycleCounterZ0Z_1 ));
    InMux I__694 (
            .O(N__3052),
            .I(N__3037));
    InMux I__693 (
            .O(N__3051),
            .I(N__3028));
    InMux I__692 (
            .O(N__3050),
            .I(N__3028));
    InMux I__691 (
            .O(N__3049),
            .I(N__3028));
    InMux I__690 (
            .O(N__3048),
            .I(N__3028));
    InMux I__689 (
            .O(N__3047),
            .I(N__3025));
    InMux I__688 (
            .O(N__3046),
            .I(N__3020));
    InMux I__687 (
            .O(N__3045),
            .I(N__3020));
    InMux I__686 (
            .O(N__3044),
            .I(N__3015));
    InMux I__685 (
            .O(N__3043),
            .I(N__3015));
    InMux I__684 (
            .O(N__3042),
            .I(N__3008));
    InMux I__683 (
            .O(N__3041),
            .I(N__3008));
    InMux I__682 (
            .O(N__3040),
            .I(N__3008));
    LocalMux I__681 (
            .O(N__3037),
            .I(N__3003));
    LocalMux I__680 (
            .O(N__3028),
            .I(N__3003));
    LocalMux I__679 (
            .O(N__3025),
            .I(uartRxInst_rState_0));
    LocalMux I__678 (
            .O(N__3020),
            .I(uartRxInst_rState_0));
    LocalMux I__677 (
            .O(N__3015),
            .I(uartRxInst_rState_0));
    LocalMux I__676 (
            .O(N__3008),
            .I(uartRxInst_rState_0));
    Odrv4 I__675 (
            .O(N__3003),
            .I(uartRxInst_rState_0));
    CascadeMux I__674 (
            .O(N__2992),
            .I(\uartRxInst.g0_0_5_cascade_ ));
    InMux I__673 (
            .O(N__2989),
            .I(N__2986));
    LocalMux I__672 (
            .O(N__2986),
            .I(\uartRxInst.g0_0_4 ));
    InMux I__671 (
            .O(N__2983),
            .I(N__2973));
    InMux I__670 (
            .O(N__2982),
            .I(N__2973));
    CascadeMux I__669 (
            .O(N__2981),
            .I(N__2969));
    InMux I__668 (
            .O(N__2980),
            .I(N__2964));
    InMux I__667 (
            .O(N__2979),
            .I(N__2964));
    InMux I__666 (
            .O(N__2978),
            .I(N__2961));
    LocalMux I__665 (
            .O(N__2973),
            .I(N__2958));
    InMux I__664 (
            .O(N__2972),
            .I(N__2953));
    InMux I__663 (
            .O(N__2969),
            .I(N__2953));
    LocalMux I__662 (
            .O(N__2964),
            .I(N__2950));
    LocalMux I__661 (
            .O(N__2961),
            .I(N__2947));
    Span4Mux_h I__660 (
            .O(N__2958),
            .I(N__2942));
    LocalMux I__659 (
            .O(N__2953),
            .I(N__2942));
    Span4Mux_v I__658 (
            .O(N__2950),
            .I(N__2939));
    Span4Mux_v I__657 (
            .O(N__2947),
            .I(N__2936));
    Span4Mux_v I__656 (
            .O(N__2942),
            .I(N__2933));
    Odrv4 I__655 (
            .O(N__2939),
            .I(i_UART_RX_c));
    Odrv4 I__654 (
            .O(N__2936),
            .I(i_UART_RX_c));
    Odrv4 I__653 (
            .O(N__2933),
            .I(i_UART_RX_c));
    CascadeMux I__652 (
            .O(N__2926),
            .I(N__2919));
    InMux I__651 (
            .O(N__2925),
            .I(N__2911));
    InMux I__650 (
            .O(N__2924),
            .I(N__2911));
    CascadeMux I__649 (
            .O(N__2923),
            .I(N__2905));
    CascadeMux I__648 (
            .O(N__2922),
            .I(N__2902));
    InMux I__647 (
            .O(N__2919),
            .I(N__2898));
    InMux I__646 (
            .O(N__2918),
            .I(N__2893));
    InMux I__645 (
            .O(N__2917),
            .I(N__2893));
    InMux I__644 (
            .O(N__2916),
            .I(N__2890));
    LocalMux I__643 (
            .O(N__2911),
            .I(N__2887));
    InMux I__642 (
            .O(N__2910),
            .I(N__2882));
    InMux I__641 (
            .O(N__2909),
            .I(N__2882));
    InMux I__640 (
            .O(N__2908),
            .I(N__2873));
    InMux I__639 (
            .O(N__2905),
            .I(N__2873));
    InMux I__638 (
            .O(N__2902),
            .I(N__2873));
    InMux I__637 (
            .O(N__2901),
            .I(N__2873));
    LocalMux I__636 (
            .O(N__2898),
            .I(uartRxInst_rState_1));
    LocalMux I__635 (
            .O(N__2893),
            .I(uartRxInst_rState_1));
    LocalMux I__634 (
            .O(N__2890),
            .I(uartRxInst_rState_1));
    Odrv4 I__633 (
            .O(N__2887),
            .I(uartRxInst_rState_1));
    LocalMux I__632 (
            .O(N__2882),
            .I(uartRxInst_rState_1));
    LocalMux I__631 (
            .O(N__2873),
            .I(uartRxInst_rState_1));
    CascadeMux I__630 (
            .O(N__2860),
            .I(\uartRxInst.N_83_0_i_0_cascade_ ));
    InMux I__629 (
            .O(N__2857),
            .I(N__2854));
    LocalMux I__628 (
            .O(N__2854),
            .I(\uartRxInst.rCycleCounter_s_3 ));
    InMux I__627 (
            .O(N__2851),
            .I(N__2842));
    InMux I__626 (
            .O(N__2850),
            .I(N__2835));
    InMux I__625 (
            .O(N__2849),
            .I(N__2835));
    InMux I__624 (
            .O(N__2848),
            .I(N__2835));
    InMux I__623 (
            .O(N__2847),
            .I(N__2828));
    InMux I__622 (
            .O(N__2846),
            .I(N__2828));
    InMux I__621 (
            .O(N__2845),
            .I(N__2828));
    LocalMux I__620 (
            .O(N__2842),
            .I(\uartRxInst.N_83_0_i_0 ));
    LocalMux I__619 (
            .O(N__2835),
            .I(\uartRxInst.N_83_0_i_0 ));
    LocalMux I__618 (
            .O(N__2828),
            .I(\uartRxInst.N_83_0_i_0 ));
    InMux I__617 (
            .O(N__2821),
            .I(N__2814));
    InMux I__616 (
            .O(N__2820),
            .I(N__2811));
    InMux I__615 (
            .O(N__2819),
            .I(N__2804));
    InMux I__614 (
            .O(N__2818),
            .I(N__2804));
    InMux I__613 (
            .O(N__2817),
            .I(N__2804));
    LocalMux I__612 (
            .O(N__2814),
            .I(\uartRxInst.rCycleCounterZ0Z_0 ));
    LocalMux I__611 (
            .O(N__2811),
            .I(\uartRxInst.rCycleCounterZ0Z_0 ));
    LocalMux I__610 (
            .O(N__2804),
            .I(\uartRxInst.rCycleCounterZ0Z_0 ));
    ClkMux I__609 (
            .O(N__2797),
            .I(N__2749));
    ClkMux I__608 (
            .O(N__2796),
            .I(N__2749));
    ClkMux I__607 (
            .O(N__2795),
            .I(N__2749));
    ClkMux I__606 (
            .O(N__2794),
            .I(N__2749));
    ClkMux I__605 (
            .O(N__2793),
            .I(N__2749));
    ClkMux I__604 (
            .O(N__2792),
            .I(N__2749));
    ClkMux I__603 (
            .O(N__2791),
            .I(N__2749));
    ClkMux I__602 (
            .O(N__2790),
            .I(N__2749));
    ClkMux I__601 (
            .O(N__2789),
            .I(N__2749));
    ClkMux I__600 (
            .O(N__2788),
            .I(N__2749));
    ClkMux I__599 (
            .O(N__2787),
            .I(N__2749));
    ClkMux I__598 (
            .O(N__2786),
            .I(N__2749));
    ClkMux I__597 (
            .O(N__2785),
            .I(N__2749));
    ClkMux I__596 (
            .O(N__2784),
            .I(N__2749));
    ClkMux I__595 (
            .O(N__2783),
            .I(N__2749));
    ClkMux I__594 (
            .O(N__2782),
            .I(N__2749));
    GlobalMux I__593 (
            .O(N__2749),
            .I(N__2746));
    gio2CtrlBuf I__592 (
            .O(N__2746),
            .I(i_Clk_c_g));
    CEMux I__591 (
            .O(N__2743),
            .I(N__2739));
    CEMux I__590 (
            .O(N__2742),
            .I(N__2736));
    LocalMux I__589 (
            .O(N__2739),
            .I(N__2732));
    LocalMux I__588 (
            .O(N__2736),
            .I(N__2729));
    CEMux I__587 (
            .O(N__2735),
            .I(N__2726));
    Span4Mux_v I__586 (
            .O(N__2732),
            .I(N__2723));
    Span4Mux_v I__585 (
            .O(N__2729),
            .I(N__2720));
    LocalMux I__584 (
            .O(N__2726),
            .I(N__2717));
    Odrv4 I__583 (
            .O(N__2723),
            .I(\uartRxInst.rCycleCountere_0_i ));
    Odrv4 I__582 (
            .O(N__2720),
            .I(\uartRxInst.rCycleCountere_0_i ));
    Odrv4 I__581 (
            .O(N__2717),
            .I(\uartRxInst.rCycleCountere_0_i ));
    InMux I__580 (
            .O(N__2710),
            .I(N__2704));
    InMux I__579 (
            .O(N__2709),
            .I(N__2701));
    InMux I__578 (
            .O(N__2708),
            .I(N__2696));
    InMux I__577 (
            .O(N__2707),
            .I(N__2696));
    LocalMux I__576 (
            .O(N__2704),
            .I(\uartRxInst.rCycleCounterZ0Z_2 ));
    LocalMux I__575 (
            .O(N__2701),
            .I(\uartRxInst.rCycleCounterZ0Z_2 ));
    LocalMux I__574 (
            .O(N__2696),
            .I(\uartRxInst.rCycleCounterZ0Z_2 ));
    CascadeMux I__573 (
            .O(N__2689),
            .I(N__2686));
    InMux I__572 (
            .O(N__2686),
            .I(N__2680));
    InMux I__571 (
            .O(N__2685),
            .I(N__2677));
    InMux I__570 (
            .O(N__2684),
            .I(N__2674));
    InMux I__569 (
            .O(N__2683),
            .I(N__2671));
    LocalMux I__568 (
            .O(N__2680),
            .I(\uartRxInst.rCycleCounterZ0Z_7 ));
    LocalMux I__567 (
            .O(N__2677),
            .I(\uartRxInst.rCycleCounterZ0Z_7 ));
    LocalMux I__566 (
            .O(N__2674),
            .I(\uartRxInst.rCycleCounterZ0Z_7 ));
    LocalMux I__565 (
            .O(N__2671),
            .I(\uartRxInst.rCycleCounterZ0Z_7 ));
    CascadeMux I__564 (
            .O(N__2662),
            .I(N__2657));
    CascadeMux I__563 (
            .O(N__2661),
            .I(N__2653));
    InMux I__562 (
            .O(N__2660),
            .I(N__2650));
    InMux I__561 (
            .O(N__2657),
            .I(N__2647));
    InMux I__560 (
            .O(N__2656),
            .I(N__2642));
    InMux I__559 (
            .O(N__2653),
            .I(N__2642));
    LocalMux I__558 (
            .O(N__2650),
            .I(\uartRxInst.rCycleCounterZ0Z_3 ));
    LocalMux I__557 (
            .O(N__2647),
            .I(\uartRxInst.rCycleCounterZ0Z_3 ));
    LocalMux I__556 (
            .O(N__2642),
            .I(\uartRxInst.rCycleCounterZ0Z_3 ));
    InMux I__555 (
            .O(N__2635),
            .I(N__2629));
    InMux I__554 (
            .O(N__2634),
            .I(N__2626));
    InMux I__553 (
            .O(N__2633),
            .I(N__2623));
    InMux I__552 (
            .O(N__2632),
            .I(N__2620));
    LocalMux I__551 (
            .O(N__2629),
            .I(\uartRxInst.rCycleCounterZ0Z_6 ));
    LocalMux I__550 (
            .O(N__2626),
            .I(\uartRxInst.rCycleCounterZ0Z_6 ));
    LocalMux I__549 (
            .O(N__2623),
            .I(\uartRxInst.rCycleCounterZ0Z_6 ));
    LocalMux I__548 (
            .O(N__2620),
            .I(\uartRxInst.rCycleCounterZ0Z_6 ));
    InMux I__547 (
            .O(N__2611),
            .I(N__2608));
    LocalMux I__546 (
            .O(N__2608),
            .I(G_11_i_a3_0_5));
    CEMux I__545 (
            .O(N__2605),
            .I(N__2602));
    LocalMux I__544 (
            .O(N__2602),
            .I(N__2599));
    Span4Mux_v I__543 (
            .O(N__2599),
            .I(N__2596));
    Odrv4 I__542 (
            .O(N__2596),
            .I(CONSTANT_ZERO_NET));
    InMux I__541 (
            .O(N__2593),
            .I(N__2590));
    LocalMux I__540 (
            .O(N__2590),
            .I(G_11_i_a3_0_6));
    CascadeMux I__539 (
            .O(N__2587),
            .I(G_11_i_a3_0_4_cascade_));
    CascadeMux I__538 (
            .O(N__2584),
            .I(N__2581));
    InMux I__537 (
            .O(N__2581),
            .I(N__2577));
    InMux I__536 (
            .O(N__2580),
            .I(N__2574));
    LocalMux I__535 (
            .O(N__2577),
            .I(uartRxInst_un1_rData_0_sqmuxa_0));
    LocalMux I__534 (
            .O(N__2574),
            .I(uartRxInst_un1_rData_0_sqmuxa_0));
    InMux I__533 (
            .O(N__2569),
            .I(N__2566));
    LocalMux I__532 (
            .O(N__2566),
            .I(N__2563));
    Odrv4 I__531 (
            .O(N__2563),
            .I(N_5));
    CEMux I__530 (
            .O(N__2560),
            .I(N__2557));
    LocalMux I__529 (
            .O(N__2557),
            .I(N__2554));
    Span4Mux_s3_h I__528 (
            .O(N__2554),
            .I(N__2551));
    Odrv4 I__527 (
            .O(N__2551),
            .I(\uartRxInst.un1_rCycleCounter_2_sqmuxa_0 ));
    CascadeMux I__526 (
            .O(N__2548),
            .I(N__2541));
    InMux I__525 (
            .O(N__2547),
            .I(N__2538));
    InMux I__524 (
            .O(N__2546),
            .I(N__2531));
    InMux I__523 (
            .O(N__2545),
            .I(N__2531));
    InMux I__522 (
            .O(N__2544),
            .I(N__2531));
    InMux I__521 (
            .O(N__2541),
            .I(N__2528));
    LocalMux I__520 (
            .O(N__2538),
            .I(\uartRxInst.rCycleCounterZ0Z_5 ));
    LocalMux I__519 (
            .O(N__2531),
            .I(\uartRxInst.rCycleCounterZ0Z_5 ));
    LocalMux I__518 (
            .O(N__2528),
            .I(\uartRxInst.rCycleCounterZ0Z_5 ));
    InMux I__517 (
            .O(N__2521),
            .I(N__2514));
    InMux I__516 (
            .O(N__2520),
            .I(N__2509));
    InMux I__515 (
            .O(N__2519),
            .I(N__2509));
    InMux I__514 (
            .O(N__2518),
            .I(N__2504));
    InMux I__513 (
            .O(N__2517),
            .I(N__2504));
    LocalMux I__512 (
            .O(N__2514),
            .I(\uartRxInst.rCycleCounterZ0Z_4 ));
    LocalMux I__511 (
            .O(N__2509),
            .I(\uartRxInst.rCycleCounterZ0Z_4 ));
    LocalMux I__510 (
            .O(N__2504),
            .I(\uartRxInst.rCycleCounterZ0Z_4 ));
    CascadeMux I__509 (
            .O(N__2497),
            .I(\uartRxInst.un12_rstate_3_cascade_ ));
    InMux I__508 (
            .O(N__2494),
            .I(N__2488));
    InMux I__507 (
            .O(N__2493),
            .I(N__2481));
    InMux I__506 (
            .O(N__2492),
            .I(N__2481));
    InMux I__505 (
            .O(N__2491),
            .I(N__2481));
    LocalMux I__504 (
            .O(N__2488),
            .I(\uartRxInst.N_83_0_i ));
    LocalMux I__503 (
            .O(N__2481),
            .I(\uartRxInst.N_83_0_i ));
    CascadeMux I__502 (
            .O(N__2476),
            .I(\uartRxInst.N_83_0_i_cascade_ ));
    InMux I__501 (
            .O(N__2473),
            .I(N__2467));
    InMux I__500 (
            .O(N__2472),
            .I(N__2467));
    LocalMux I__499 (
            .O(N__2467),
            .I(\uartRxInst.rState_0_sqmuxa_1_1 ));
    CascadeMux I__498 (
            .O(N__2464),
            .I(N__2460));
    InMux I__497 (
            .O(N__2463),
            .I(N__2452));
    InMux I__496 (
            .O(N__2460),
            .I(N__2452));
    InMux I__495 (
            .O(N__2459),
            .I(N__2452));
    LocalMux I__494 (
            .O(N__2452),
            .I(\uartRxInst.rDataCounter_0_sqmuxa ));
    InMux I__493 (
            .O(N__2449),
            .I(N__2446));
    LocalMux I__492 (
            .O(N__2446),
            .I(\uartRxInst.rCycleCounter_cry_0_THRU_CO ));
    SRMux I__491 (
            .O(N__2443),
            .I(N__2439));
    InMux I__490 (
            .O(N__2442),
            .I(N__2436));
    LocalMux I__489 (
            .O(N__2439),
            .I(N__2433));
    LocalMux I__488 (
            .O(N__2436),
            .I(N__2430));
    Odrv12 I__487 (
            .O(N__2433),
            .I(\uartRxInst.rstateZ0 ));
    Odrv4 I__486 (
            .O(N__2430),
            .I(\uartRxInst.rstateZ0 ));
    InMux I__485 (
            .O(N__2425),
            .I(N__2422));
    LocalMux I__484 (
            .O(N__2422),
            .I(\uartRxInst.rCycleCounter_s_2 ));
    CascadeMux I__483 (
            .O(N__2419),
            .I(pEcho_rRamAddress_2_5_cascade_));
    CascadeMux I__482 (
            .O(N__2416),
            .I(N__2413));
    InMux I__481 (
            .O(N__2413),
            .I(N__2409));
    InMux I__480 (
            .O(N__2412),
            .I(N__2406));
    LocalMux I__479 (
            .O(N__2409),
            .I(rRamAddressZ0Z_5));
    LocalMux I__478 (
            .O(N__2406),
            .I(rRamAddressZ0Z_5));
    CascadeMux I__477 (
            .O(N__2401),
            .I(N__2398));
    InMux I__476 (
            .O(N__2398),
            .I(N__2394));
    InMux I__475 (
            .O(N__2397),
            .I(N__2391));
    LocalMux I__474 (
            .O(N__2394),
            .I(pEcho_rRamAddress_2_3));
    LocalMux I__473 (
            .O(N__2391),
            .I(pEcho_rRamAddress_2_3));
    CascadeMux I__472 (
            .O(N__2386),
            .I(N__2383));
    InMux I__471 (
            .O(N__2383),
            .I(N__2379));
    InMux I__470 (
            .O(N__2382),
            .I(N__2376));
    LocalMux I__469 (
            .O(N__2379),
            .I(rRamAddressZ0Z_3));
    LocalMux I__468 (
            .O(N__2376),
            .I(rRamAddressZ0Z_3));
    InMux I__467 (
            .O(N__2371),
            .I(N__2368));
    LocalMux I__466 (
            .O(N__2368),
            .I(rRamReadData_0));
    CascadeMux I__465 (
            .O(N__2365),
            .I(N__2362));
    InMux I__464 (
            .O(N__2362),
            .I(N__2359));
    LocalMux I__463 (
            .O(N__2359),
            .I(N__2356));
    Odrv4 I__462 (
            .O(N__2356),
            .I(rTxByteZ0Z_4));
    InMux I__461 (
            .O(N__2353),
            .I(N__2350));
    LocalMux I__460 (
            .O(N__2350),
            .I(rRamReadData_1));
    InMux I__459 (
            .O(N__2347),
            .I(N__2344));
    LocalMux I__458 (
            .O(N__2344),
            .I(rTxByteZ0Z_5));
    InMux I__457 (
            .O(N__2341),
            .I(N__2338));
    LocalMux I__456 (
            .O(N__2338),
            .I(rRamReadData_2));
    CascadeMux I__455 (
            .O(N__2335),
            .I(N__2332));
    InMux I__454 (
            .O(N__2332),
            .I(N__2329));
    LocalMux I__453 (
            .O(N__2329),
            .I(N__2326));
    Odrv4 I__452 (
            .O(N__2326),
            .I(rTxByteZ0Z_6));
    InMux I__451 (
            .O(N__2323),
            .I(N__2320));
    LocalMux I__450 (
            .O(N__2320),
            .I(rRamReadData_3));
    CascadeMux I__449 (
            .O(N__2317),
            .I(N__2314));
    InMux I__448 (
            .O(N__2314),
            .I(N__2311));
    LocalMux I__447 (
            .O(N__2311),
            .I(N__2308));
    Odrv4 I__446 (
            .O(N__2308),
            .I(rTxByteZ0Z_7));
    CEMux I__445 (
            .O(N__2305),
            .I(N__2301));
    CascadeMux I__444 (
            .O(N__2304),
            .I(N__2294));
    LocalMux I__443 (
            .O(N__2301),
            .I(N__2291));
    InMux I__442 (
            .O(N__2300),
            .I(N__2288));
    InMux I__441 (
            .O(N__2299),
            .I(N__2285));
    InMux I__440 (
            .O(N__2298),
            .I(N__2282));
    InMux I__439 (
            .O(N__2297),
            .I(N__2279));
    InMux I__438 (
            .O(N__2294),
            .I(N__2276));
    Odrv4 I__437 (
            .O(N__2291),
            .I(rRxReady));
    LocalMux I__436 (
            .O(N__2288),
            .I(rRxReady));
    LocalMux I__435 (
            .O(N__2285),
            .I(rRxReady));
    LocalMux I__434 (
            .O(N__2282),
            .I(rRxReady));
    LocalMux I__433 (
            .O(N__2279),
            .I(rRxReady));
    LocalMux I__432 (
            .O(N__2276),
            .I(rRxReady));
    InMux I__431 (
            .O(N__2263),
            .I(\uartRxInst.rCycleCounter_cry_6 ));
    CascadeMux I__430 (
            .O(N__2260),
            .I(N__2257));
    InMux I__429 (
            .O(N__2257),
            .I(N__2254));
    LocalMux I__428 (
            .O(N__2254),
            .I(N__2249));
    InMux I__427 (
            .O(N__2253),
            .I(N__2246));
    InMux I__426 (
            .O(N__2252),
            .I(N__2243));
    Odrv4 I__425 (
            .O(N__2249),
            .I(rRamAddressZ0Z_0));
    LocalMux I__424 (
            .O(N__2246),
            .I(rRamAddressZ0Z_0));
    LocalMux I__423 (
            .O(N__2243),
            .I(rRamAddressZ0Z_0));
    CascadeMux I__422 (
            .O(N__2236),
            .I(N__2233));
    InMux I__421 (
            .O(N__2233),
            .I(N__2230));
    LocalMux I__420 (
            .O(N__2230),
            .I(pEcho_rRamAddress_2_0));
    CascadeMux I__419 (
            .O(N__2227),
            .I(N__2224));
    InMux I__418 (
            .O(N__2224),
            .I(N__2221));
    LocalMux I__417 (
            .O(N__2221),
            .I(N__2217));
    InMux I__416 (
            .O(N__2220),
            .I(N__2214));
    Odrv4 I__415 (
            .O(N__2217),
            .I(rRamAddressZ0Z_1));
    LocalMux I__414 (
            .O(N__2214),
            .I(rRamAddressZ0Z_1));
    CascadeMux I__413 (
            .O(N__2209),
            .I(N__2206));
    InMux I__412 (
            .O(N__2206),
            .I(N__2202));
    InMux I__411 (
            .O(N__2205),
            .I(N__2199));
    LocalMux I__410 (
            .O(N__2202),
            .I(pEcho_rRamAddress_2_1));
    LocalMux I__409 (
            .O(N__2199),
            .I(pEcho_rRamAddress_2_1));
    InMux I__408 (
            .O(N__2194),
            .I(pEcho_rRamAddress_2_cry_0));
    CascadeMux I__407 (
            .O(N__2191),
            .I(N__2188));
    InMux I__406 (
            .O(N__2188),
            .I(N__2185));
    LocalMux I__405 (
            .O(N__2185),
            .I(N__2181));
    InMux I__404 (
            .O(N__2184),
            .I(N__2178));
    Odrv4 I__403 (
            .O(N__2181),
            .I(rRamAddressZ0Z_2));
    LocalMux I__402 (
            .O(N__2178),
            .I(rRamAddressZ0Z_2));
    CascadeMux I__401 (
            .O(N__2173),
            .I(N__2170));
    InMux I__400 (
            .O(N__2170),
            .I(N__2166));
    InMux I__399 (
            .O(N__2169),
            .I(N__2163));
    LocalMux I__398 (
            .O(N__2166),
            .I(pEcho_rRamAddress_2_2));
    LocalMux I__397 (
            .O(N__2163),
            .I(pEcho_rRamAddress_2_2));
    InMux I__396 (
            .O(N__2158),
            .I(pEcho_rRamAddress_2_cry_1));
    InMux I__395 (
            .O(N__2155),
            .I(pEcho_rRamAddress_2_cry_2));
    CascadeMux I__394 (
            .O(N__2152),
            .I(N__2149));
    InMux I__393 (
            .O(N__2149),
            .I(N__2146));
    LocalMux I__392 (
            .O(N__2146),
            .I(N__2142));
    InMux I__391 (
            .O(N__2145),
            .I(N__2139));
    Odrv4 I__390 (
            .O(N__2142),
            .I(rRamAddressZ0Z_4));
    LocalMux I__389 (
            .O(N__2139),
            .I(rRamAddressZ0Z_4));
    CascadeMux I__388 (
            .O(N__2134),
            .I(N__2131));
    InMux I__387 (
            .O(N__2131),
            .I(N__2127));
    InMux I__386 (
            .O(N__2130),
            .I(N__2124));
    LocalMux I__385 (
            .O(N__2127),
            .I(pEcho_rRamAddress_2_4));
    LocalMux I__384 (
            .O(N__2124),
            .I(pEcho_rRamAddress_2_4));
    InMux I__383 (
            .O(N__2119),
            .I(pEcho_rRamAddress_2_cry_3));
    InMux I__382 (
            .O(N__2116),
            .I(pEcho_rRamAddress_2_cry_4));
    CascadeMux I__381 (
            .O(N__2113),
            .I(N__2110));
    InMux I__380 (
            .O(N__2110),
            .I(N__2107));
    LocalMux I__379 (
            .O(N__2107),
            .I(pEcho_rRamAddress_2_5));
    CascadeMux I__378 (
            .O(N__2104),
            .I(N__2100));
    InMux I__377 (
            .O(N__2103),
            .I(N__2096));
    InMux I__376 (
            .O(N__2100),
            .I(N__2091));
    InMux I__375 (
            .O(N__2099),
            .I(N__2091));
    LocalMux I__374 (
            .O(N__2096),
            .I(\uartRxInst.rDataCounterZ0Z_1 ));
    LocalMux I__373 (
            .O(N__2091),
            .I(\uartRxInst.rDataCounterZ0Z_1 ));
    InMux I__372 (
            .O(N__2086),
            .I(N__2083));
    LocalMux I__371 (
            .O(N__2083),
            .I(N__2077));
    InMux I__370 (
            .O(N__2082),
            .I(N__2070));
    InMux I__369 (
            .O(N__2081),
            .I(N__2070));
    InMux I__368 (
            .O(N__2080),
            .I(N__2070));
    Odrv4 I__367 (
            .O(N__2077),
            .I(\uartRxInst.rDataCounterZ0Z_0 ));
    LocalMux I__366 (
            .O(N__2070),
            .I(\uartRxInst.rDataCounterZ0Z_0 ));
    InMux I__365 (
            .O(N__2065),
            .I(N__2062));
    LocalMux I__364 (
            .O(N__2062),
            .I(\uartRxInst.CO1_0 ));
    InMux I__363 (
            .O(N__2059),
            .I(\uartRxInst.rCycleCounter_cry_0 ));
    InMux I__362 (
            .O(N__2056),
            .I(\uartRxInst.rCycleCounter_cry_1 ));
    InMux I__361 (
            .O(N__2053),
            .I(\uartRxInst.rCycleCounter_cry_2 ));
    InMux I__360 (
            .O(N__2050),
            .I(N__2047));
    LocalMux I__359 (
            .O(N__2047),
            .I(\uartRxInst.rCycleCounter_cry_3_THRU_CO ));
    InMux I__358 (
            .O(N__2044),
            .I(\uartRxInst.rCycleCounter_cry_3 ));
    InMux I__357 (
            .O(N__2041),
            .I(N__2038));
    LocalMux I__356 (
            .O(N__2038),
            .I(\uartRxInst.rCycleCounter_s_5 ));
    InMux I__355 (
            .O(N__2035),
            .I(\uartRxInst.rCycleCounter_cry_4 ));
    CascadeMux I__354 (
            .O(N__2032),
            .I(N__2027));
    CascadeMux I__353 (
            .O(N__2031),
            .I(N__2024));
    CascadeMux I__352 (
            .O(N__2030),
            .I(N__2021));
    InMux I__351 (
            .O(N__2027),
            .I(N__2011));
    InMux I__350 (
            .O(N__2024),
            .I(N__2011));
    InMux I__349 (
            .O(N__2021),
            .I(N__2011));
    CascadeMux I__348 (
            .O(N__2020),
            .I(N__2006));
    CascadeMux I__347 (
            .O(N__2019),
            .I(N__2003));
    CascadeMux I__346 (
            .O(N__2018),
            .I(N__2000));
    LocalMux I__345 (
            .O(N__2011),
            .I(N__1997));
    SRMux I__344 (
            .O(N__2010),
            .I(N__1994));
    SRMux I__343 (
            .O(N__2009),
            .I(N__1991));
    InMux I__342 (
            .O(N__2006),
            .I(N__1984));
    InMux I__341 (
            .O(N__2003),
            .I(N__1984));
    InMux I__340 (
            .O(N__2000),
            .I(N__1984));
    Span4Mux_v I__339 (
            .O(N__1997),
            .I(N__1979));
    LocalMux I__338 (
            .O(N__1994),
            .I(N__1979));
    LocalMux I__337 (
            .O(N__1991),
            .I(N__1976));
    LocalMux I__336 (
            .O(N__1984),
            .I(N__1973));
    Span4Mux_h I__335 (
            .O(N__1979),
            .I(N__1970));
    Span4Mux_v I__334 (
            .O(N__1976),
            .I(N__1967));
    Odrv12 I__333 (
            .O(N__1973),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__332 (
            .O(N__1970),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__331 (
            .O(N__1967),
            .I(CONSTANT_ONE_NET));
    InMux I__330 (
            .O(N__1960),
            .I(N__1957));
    LocalMux I__329 (
            .O(N__1957),
            .I(\uartRxInst.rCycleCounter_s_6 ));
    InMux I__328 (
            .O(N__1954),
            .I(\uartRxInst.rCycleCounter_cry_5 ));
    InMux I__327 (
            .O(N__1951),
            .I(N__1943));
    InMux I__326 (
            .O(N__1950),
            .I(N__1943));
    InMux I__325 (
            .O(N__1949),
            .I(N__1940));
    InMux I__324 (
            .O(N__1948),
            .I(N__1937));
    LocalMux I__323 (
            .O(N__1943),
            .I(\uartTxInst.rBitIndexZ0Z_1 ));
    LocalMux I__322 (
            .O(N__1940),
            .I(\uartTxInst.rBitIndexZ0Z_1 ));
    LocalMux I__321 (
            .O(N__1937),
            .I(\uartTxInst.rBitIndexZ0Z_1 ));
    CascadeMux I__320 (
            .O(N__1930),
            .I(N__1926));
    InMux I__319 (
            .O(N__1929),
            .I(N__1923));
    InMux I__318 (
            .O(N__1926),
            .I(N__1920));
    LocalMux I__317 (
            .O(N__1923),
            .I(\uartTxInst.rTxByte_0_4 ));
    LocalMux I__316 (
            .O(N__1920),
            .I(\uartTxInst.rTxByte_0_4 ));
    InMux I__315 (
            .O(N__1915),
            .I(N__1911));
    InMux I__314 (
            .O(N__1914),
            .I(N__1908));
    LocalMux I__313 (
            .O(N__1911),
            .I(\uartTxInst.rTxByte_0_6 ));
    LocalMux I__312 (
            .O(N__1908),
            .I(\uartTxInst.rTxByte_0_6 ));
    InMux I__311 (
            .O(N__1903),
            .I(N__1896));
    InMux I__310 (
            .O(N__1902),
            .I(N__1893));
    InMux I__309 (
            .O(N__1901),
            .I(N__1890));
    InMux I__308 (
            .O(N__1900),
            .I(N__1885));
    InMux I__307 (
            .O(N__1899),
            .I(N__1885));
    LocalMux I__306 (
            .O(N__1896),
            .I(N__1882));
    LocalMux I__305 (
            .O(N__1893),
            .I(\uartTxInst.rBitIndexZ1Z_0 ));
    LocalMux I__304 (
            .O(N__1890),
            .I(\uartTxInst.rBitIndexZ1Z_0 ));
    LocalMux I__303 (
            .O(N__1885),
            .I(\uartTxInst.rBitIndexZ1Z_0 ));
    Odrv4 I__302 (
            .O(N__1882),
            .I(\uartTxInst.rBitIndexZ1Z_0 ));
    InMux I__301 (
            .O(N__1873),
            .I(N__1869));
    InMux I__300 (
            .O(N__1872),
            .I(N__1866));
    LocalMux I__299 (
            .O(N__1869),
            .I(\uartTxInst.rTxByte_0_7 ));
    LocalMux I__298 (
            .O(N__1866),
            .I(\uartTxInst.rTxByte_0_7 ));
    CascadeMux I__297 (
            .O(N__1861),
            .I(\uartTxInst.oSerial_3_6_i_m2_ns_1_cascade_ ));
    CascadeMux I__296 (
            .O(N__1858),
            .I(N__1855));
    InMux I__295 (
            .O(N__1855),
            .I(N__1851));
    InMux I__294 (
            .O(N__1854),
            .I(N__1848));
    LocalMux I__293 (
            .O(N__1851),
            .I(\uartTxInst.rTxByte_0_5 ));
    LocalMux I__292 (
            .O(N__1848),
            .I(\uartTxInst.rTxByte_0_5 ));
    InMux I__291 (
            .O(N__1843),
            .I(N__1838));
    InMux I__290 (
            .O(N__1842),
            .I(N__1835));
    InMux I__289 (
            .O(N__1841),
            .I(N__1832));
    LocalMux I__288 (
            .O(N__1838),
            .I(\uartTxInst.rBitIndexZ0Z_2 ));
    LocalMux I__287 (
            .O(N__1835),
            .I(\uartTxInst.rBitIndexZ0Z_2 ));
    LocalMux I__286 (
            .O(N__1832),
            .I(\uartTxInst.rBitIndexZ0Z_2 ));
    CascadeMux I__285 (
            .O(N__1825),
            .I(\uartTxInst.N_35_cascade_ ));
    InMux I__284 (
            .O(N__1822),
            .I(N__1812));
    InMux I__283 (
            .O(N__1821),
            .I(N__1809));
    InMux I__282 (
            .O(N__1820),
            .I(N__1806));
    InMux I__281 (
            .O(N__1819),
            .I(N__1797));
    InMux I__280 (
            .O(N__1818),
            .I(N__1797));
    InMux I__279 (
            .O(N__1817),
            .I(N__1797));
    InMux I__278 (
            .O(N__1816),
            .I(N__1797));
    InMux I__277 (
            .O(N__1815),
            .I(N__1794));
    LocalMux I__276 (
            .O(N__1812),
            .I(\uartTxInst.rTxStateZ0Z_0 ));
    LocalMux I__275 (
            .O(N__1809),
            .I(\uartTxInst.rTxStateZ0Z_0 ));
    LocalMux I__274 (
            .O(N__1806),
            .I(\uartTxInst.rTxStateZ0Z_0 ));
    LocalMux I__273 (
            .O(N__1797),
            .I(\uartTxInst.rTxStateZ0Z_0 ));
    LocalMux I__272 (
            .O(N__1794),
            .I(\uartTxInst.rTxStateZ0Z_0 ));
    InMux I__271 (
            .O(N__1783),
            .I(N__1780));
    LocalMux I__270 (
            .O(N__1780),
            .I(\uartTxInst.N_48 ));
    CascadeMux I__269 (
            .O(N__1777),
            .I(N__1774));
    InMux I__268 (
            .O(N__1774),
            .I(N__1768));
    InMux I__267 (
            .O(N__1773),
            .I(N__1768));
    LocalMux I__266 (
            .O(N__1768),
            .I(\uartRxInst.rDataCounterZ0Z_2 ));
    CascadeMux I__265 (
            .O(N__1765),
            .I(\uartRxInst.rstateZ0_cascade_ ));
    InMux I__264 (
            .O(N__1762),
            .I(N__1759));
    LocalMux I__263 (
            .O(N__1759),
            .I(\uartTxInst.N_31 ));
    CascadeMux I__262 (
            .O(N__1756),
            .I(N__1751));
    CascadeMux I__261 (
            .O(N__1755),
            .I(N__1746));
    CascadeMux I__260 (
            .O(N__1754),
            .I(N__1743));
    InMux I__259 (
            .O(N__1751),
            .I(N__1734));
    InMux I__258 (
            .O(N__1750),
            .I(N__1734));
    InMux I__257 (
            .O(N__1749),
            .I(N__1731));
    InMux I__256 (
            .O(N__1746),
            .I(N__1722));
    InMux I__255 (
            .O(N__1743),
            .I(N__1722));
    InMux I__254 (
            .O(N__1742),
            .I(N__1722));
    InMux I__253 (
            .O(N__1741),
            .I(N__1722));
    InMux I__252 (
            .O(N__1740),
            .I(N__1717));
    InMux I__251 (
            .O(N__1739),
            .I(N__1717));
    LocalMux I__250 (
            .O(N__1734),
            .I(\uartTxInst.rTxStateZ0Z_1 ));
    LocalMux I__249 (
            .O(N__1731),
            .I(\uartTxInst.rTxStateZ0Z_1 ));
    LocalMux I__248 (
            .O(N__1722),
            .I(\uartTxInst.rTxStateZ0Z_1 ));
    LocalMux I__247 (
            .O(N__1717),
            .I(\uartTxInst.rTxStateZ0Z_1 ));
    InMux I__246 (
            .O(N__1708),
            .I(N__1705));
    LocalMux I__245 (
            .O(N__1705),
            .I(\uartTxInst.un2_rclkcount_4 ));
    CascadeMux I__244 (
            .O(N__1702),
            .I(\uartTxInst.N_31_cascade_ ));
    InMux I__243 (
            .O(N__1699),
            .I(N__1696));
    LocalMux I__242 (
            .O(N__1696),
            .I(\uartTxInst.rTxState_10_0_x2_0_o2_1_1_1 ));
    CascadeMux I__241 (
            .O(N__1693),
            .I(\uartTxInst.rTxState_10_0_x2_0_o2_1_1_1_cascade_ ));
    InMux I__240 (
            .O(N__1690),
            .I(N__1686));
    InMux I__239 (
            .O(N__1689),
            .I(N__1683));
    LocalMux I__238 (
            .O(N__1686),
            .I(\uartTxInst.rTxState_10_0_x2_0_o2_d_0_1 ));
    LocalMux I__237 (
            .O(N__1683),
            .I(\uartTxInst.rTxState_10_0_x2_0_o2_d_0_1 ));
    SRMux I__236 (
            .O(N__1678),
            .I(N__1673));
    CascadeMux I__235 (
            .O(N__1677),
            .I(N__1662));
    CascadeMux I__234 (
            .O(N__1676),
            .I(N__1657));
    LocalMux I__233 (
            .O(N__1673),
            .I(N__1653));
    InMux I__232 (
            .O(N__1672),
            .I(N__1650));
    InMux I__231 (
            .O(N__1671),
            .I(N__1639));
    InMux I__230 (
            .O(N__1670),
            .I(N__1639));
    InMux I__229 (
            .O(N__1669),
            .I(N__1639));
    InMux I__228 (
            .O(N__1668),
            .I(N__1639));
    InMux I__227 (
            .O(N__1667),
            .I(N__1639));
    InMux I__226 (
            .O(N__1666),
            .I(N__1632));
    InMux I__225 (
            .O(N__1665),
            .I(N__1632));
    InMux I__224 (
            .O(N__1662),
            .I(N__1632));
    InMux I__223 (
            .O(N__1661),
            .I(N__1627));
    InMux I__222 (
            .O(N__1660),
            .I(N__1627));
    InMux I__221 (
            .O(N__1657),
            .I(N__1622));
    InMux I__220 (
            .O(N__1656),
            .I(N__1622));
    Odrv12 I__219 (
            .O(N__1653),
            .I(\uartTxInst.rbitindex15 ));
    LocalMux I__218 (
            .O(N__1650),
            .I(\uartTxInst.rbitindex15 ));
    LocalMux I__217 (
            .O(N__1639),
            .I(\uartTxInst.rbitindex15 ));
    LocalMux I__216 (
            .O(N__1632),
            .I(\uartTxInst.rbitindex15 ));
    LocalMux I__215 (
            .O(N__1627),
            .I(\uartTxInst.rbitindex15 ));
    LocalMux I__214 (
            .O(N__1622),
            .I(\uartTxInst.rbitindex15 ));
    InMux I__213 (
            .O(N__1609),
            .I(N__1602));
    InMux I__212 (
            .O(N__1608),
            .I(N__1593));
    InMux I__211 (
            .O(N__1607),
            .I(N__1593));
    InMux I__210 (
            .O(N__1606),
            .I(N__1593));
    InMux I__209 (
            .O(N__1605),
            .I(N__1593));
    LocalMux I__208 (
            .O(N__1602),
            .I(N__1590));
    LocalMux I__207 (
            .O(N__1593),
            .I(rTxDVZ0));
    Odrv4 I__206 (
            .O(N__1590),
            .I(rTxDVZ0));
    CascadeMux I__205 (
            .O(N__1585),
            .I(\uartRxInst.rDataCounter_RNO_0Z0Z_1_cascade_ ));
    CascadeMux I__204 (
            .O(N__1582),
            .I(\uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_ ));
    InMux I__203 (
            .O(N__1579),
            .I(N__1574));
    InMux I__202 (
            .O(N__1578),
            .I(N__1571));
    InMux I__201 (
            .O(N__1577),
            .I(N__1568));
    LocalMux I__200 (
            .O(N__1574),
            .I(\uartTxInst.rClkCountZ0Z_6 ));
    LocalMux I__199 (
            .O(N__1571),
            .I(\uartTxInst.rClkCountZ0Z_6 ));
    LocalMux I__198 (
            .O(N__1568),
            .I(\uartTxInst.rClkCountZ0Z_6 ));
    CascadeMux I__197 (
            .O(N__1561),
            .I(N__1557));
    InMux I__196 (
            .O(N__1560),
            .I(N__1552));
    InMux I__195 (
            .O(N__1557),
            .I(N__1547));
    InMux I__194 (
            .O(N__1556),
            .I(N__1547));
    InMux I__193 (
            .O(N__1555),
            .I(N__1544));
    LocalMux I__192 (
            .O(N__1552),
            .I(\uartTxInst.rClkCountZ0Z_5 ));
    LocalMux I__191 (
            .O(N__1547),
            .I(\uartTxInst.rClkCountZ0Z_5 ));
    LocalMux I__190 (
            .O(N__1544),
            .I(\uartTxInst.rClkCountZ0Z_5 ));
    CascadeMux I__189 (
            .O(N__1537),
            .I(N__1532));
    InMux I__188 (
            .O(N__1536),
            .I(N__1525));
    InMux I__187 (
            .O(N__1535),
            .I(N__1525));
    InMux I__186 (
            .O(N__1532),
            .I(N__1525));
    LocalMux I__185 (
            .O(N__1525),
            .I(\uartTxInst.un5_rclkcount_c4 ));
    InMux I__184 (
            .O(N__1522),
            .I(N__1508));
    InMux I__183 (
            .O(N__1521),
            .I(N__1508));
    InMux I__182 (
            .O(N__1520),
            .I(N__1505));
    InMux I__181 (
            .O(N__1519),
            .I(N__1500));
    InMux I__180 (
            .O(N__1518),
            .I(N__1500));
    InMux I__179 (
            .O(N__1517),
            .I(N__1497));
    InMux I__178 (
            .O(N__1516),
            .I(N__1494));
    InMux I__177 (
            .O(N__1515),
            .I(N__1487));
    InMux I__176 (
            .O(N__1514),
            .I(N__1487));
    InMux I__175 (
            .O(N__1513),
            .I(N__1487));
    LocalMux I__174 (
            .O(N__1508),
            .I(N__1484));
    LocalMux I__173 (
            .O(N__1505),
            .I(\uartTxInst.SUM_N_3_mux ));
    LocalMux I__172 (
            .O(N__1500),
            .I(\uartTxInst.SUM_N_3_mux ));
    LocalMux I__171 (
            .O(N__1497),
            .I(\uartTxInst.SUM_N_3_mux ));
    LocalMux I__170 (
            .O(N__1494),
            .I(\uartTxInst.SUM_N_3_mux ));
    LocalMux I__169 (
            .O(N__1487),
            .I(\uartTxInst.SUM_N_3_mux ));
    Odrv4 I__168 (
            .O(N__1484),
            .I(\uartTxInst.SUM_N_3_mux ));
    CascadeMux I__167 (
            .O(N__1471),
            .I(N__1468));
    InMux I__166 (
            .O(N__1468),
            .I(N__1461));
    InMux I__165 (
            .O(N__1467),
            .I(N__1458));
    InMux I__164 (
            .O(N__1466),
            .I(N__1451));
    InMux I__163 (
            .O(N__1465),
            .I(N__1451));
    InMux I__162 (
            .O(N__1464),
            .I(N__1451));
    LocalMux I__161 (
            .O(N__1461),
            .I(N__1448));
    LocalMux I__160 (
            .O(N__1458),
            .I(\uartTxInst.rClkCountZ0Z_4 ));
    LocalMux I__159 (
            .O(N__1451),
            .I(\uartTxInst.rClkCountZ0Z_4 ));
    Odrv4 I__158 (
            .O(N__1448),
            .I(\uartTxInst.rClkCountZ0Z_4 ));
    CascadeMux I__157 (
            .O(N__1441),
            .I(\uartTxInst.g2_0_cascade_ ));
    CascadeMux I__156 (
            .O(N__1438),
            .I(\uartTxInst.rBitIndex_RNO_0Z0Z_1_cascade_ ));
    InMux I__155 (
            .O(N__1435),
            .I(N__1432));
    LocalMux I__154 (
            .O(N__1432),
            .I(\uartTxInst.rTxByte_0_sqmuxa ));
    CascadeMux I__153 (
            .O(N__1429),
            .I(\uartTxInst.rTxState_10_0_i_a2_1_2_0_cascade_ ));
    IoInMux I__152 (
            .O(N__1426),
            .I(N__1423));
    LocalMux I__151 (
            .O(N__1423),
            .I(N__1420));
    IoSpan4Mux I__150 (
            .O(N__1420),
            .I(N__1416));
    CascadeMux I__149 (
            .O(N__1419),
            .I(N__1413));
    Span4Mux_s2_h I__148 (
            .O(N__1416),
            .I(N__1410));
    InMux I__147 (
            .O(N__1413),
            .I(N__1407));
    Odrv4 I__146 (
            .O(N__1410),
            .I(o_UART_TX_c));
    LocalMux I__145 (
            .O(N__1407),
            .I(o_UART_TX_c));
    CascadeMux I__144 (
            .O(N__1402),
            .I(\uartTxInst.rbitindex15_cascade_ ));
    InMux I__143 (
            .O(N__1399),
            .I(N__1388));
    InMux I__142 (
            .O(N__1398),
            .I(N__1388));
    InMux I__141 (
            .O(N__1397),
            .I(N__1388));
    InMux I__140 (
            .O(N__1396),
            .I(N__1383));
    InMux I__139 (
            .O(N__1395),
            .I(N__1383));
    LocalMux I__138 (
            .O(N__1388),
            .I(\uartTxInst.rClkCountZ0Z_1 ));
    LocalMux I__137 (
            .O(N__1383),
            .I(\uartTxInst.rClkCountZ0Z_1 ));
    CascadeMux I__136 (
            .O(N__1378),
            .I(\uartTxInst.un2_rclkcount_5_0_cascade_ ));
    InMux I__135 (
            .O(N__1375),
            .I(N__1371));
    InMux I__134 (
            .O(N__1374),
            .I(N__1368));
    LocalMux I__133 (
            .O(N__1371),
            .I(\uartTxInst.rClkCountZ0Z_7 ));
    LocalMux I__132 (
            .O(N__1368),
            .I(\uartTxInst.rClkCountZ0Z_7 ));
    InMux I__131 (
            .O(N__1363),
            .I(N__1356));
    InMux I__130 (
            .O(N__1362),
            .I(N__1356));
    InMux I__129 (
            .O(N__1361),
            .I(N__1353));
    LocalMux I__128 (
            .O(N__1356),
            .I(\uartTxInst.rClkCountZ0Z_3 ));
    LocalMux I__127 (
            .O(N__1353),
            .I(\uartTxInst.rClkCountZ0Z_3 ));
    CascadeMux I__126 (
            .O(N__1348),
            .I(N__1343));
    CascadeMux I__125 (
            .O(N__1347),
            .I(N__1340));
    InMux I__124 (
            .O(N__1346),
            .I(N__1331));
    InMux I__123 (
            .O(N__1343),
            .I(N__1331));
    InMux I__122 (
            .O(N__1340),
            .I(N__1331));
    InMux I__121 (
            .O(N__1339),
            .I(N__1326));
    InMux I__120 (
            .O(N__1338),
            .I(N__1326));
    LocalMux I__119 (
            .O(N__1331),
            .I(\uartTxInst.rClkCountZ0Z_2 ));
    LocalMux I__118 (
            .O(N__1326),
            .I(\uartTxInst.rClkCountZ0Z_2 ));
    InMux I__117 (
            .O(N__1321),
            .I(N__1306));
    InMux I__116 (
            .O(N__1320),
            .I(N__1306));
    InMux I__115 (
            .O(N__1319),
            .I(N__1306));
    InMux I__114 (
            .O(N__1318),
            .I(N__1306));
    InMux I__113 (
            .O(N__1317),
            .I(N__1299));
    InMux I__112 (
            .O(N__1316),
            .I(N__1299));
    InMux I__111 (
            .O(N__1315),
            .I(N__1299));
    LocalMux I__110 (
            .O(N__1306),
            .I(\uartTxInst.rClkCountZ0Z_0 ));
    LocalMux I__109 (
            .O(N__1299),
            .I(\uartTxInst.rClkCountZ0Z_0 ));
    CascadeMux I__108 (
            .O(N__1294),
            .I(\uartTxInst.un2_rclkcount_4_cascade_ ));
    InMux I__107 (
            .O(N__1291),
            .I(N__1288));
    LocalMux I__106 (
            .O(N__1288),
            .I(\uartTxInst.un2_rclkcount_5_0 ));
    CascadeMux I__105 (
            .O(N__1285),
            .I(\uartTxInst.un5_rclkcount_c4_cascade_ ));
    CascadeMux I__104 (
            .O(N__1282),
            .I(\uartTxInst.un5_rclkcount_ac0_11_cascade_ ));
    CascadeMux I__103 (
            .O(N__1279),
            .I(\uartTxInst.un5_rclkcount_c3_cascade_ ));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uartTxInst.rClkCount_RNIA4KC_3_LC_7_9_0 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_RNIA4KC_3_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rClkCount_RNIA4KC_3_LC_7_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uartTxInst.rClkCount_RNIA4KC_3_LC_7_9_0  (
            .in0(N__1318),
            .in1(N__1397),
            .in2(N__1347),
            .in3(N__1362),
            .lcout(\uartTxInst.un5_rclkcount_c4 ),
            .ltout(\uartTxInst.un5_rclkcount_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_RNO_0_7_LC_7_9_1 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_RNO_0_7_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rClkCount_RNO_0_7_LC_7_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uartTxInst.rClkCount_RNO_0_7_LC_7_9_1  (
            .in0(N__1579),
            .in1(N__1560),
            .in2(N__1285),
            .in3(N__1467),
            .lcout(),
            .ltout(\uartTxInst.un5_rclkcount_ac0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_7_LC_7_9_2 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_7_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rClkCount_7_LC_7_9_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \uartTxInst.rClkCount_7_LC_7_9_2  (
            .in0(N__1661),
            .in1(N__1375),
            .in2(N__1282),
            .in3(N__1519),
            .lcout(\uartTxInst.rClkCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2782),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_2_LC_7_9_3 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_2_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rClkCount_2_LC_7_9_3 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \uartTxInst.rClkCount_2_LC_7_9_3  (
            .in0(N__1399),
            .in1(N__1346),
            .in2(N__1676),
            .in3(N__1320),
            .lcout(\uartTxInst.rClkCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2782),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_RNO_0_3_LC_7_9_4 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_RNO_0_3_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rClkCount_RNO_0_3_LC_7_9_4 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \uartTxInst.rClkCount_RNO_0_3_LC_7_9_4  (
            .in0(N__1319),
            .in1(N__1398),
            .in2(N__1348),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\uartTxInst.un5_rclkcount_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_3_LC_7_9_5 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_3_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rClkCount_3_LC_7_9_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \uartTxInst.rClkCount_3_LC_7_9_5  (
            .in0(N__1363),
            .in1(N__1660),
            .in2(N__1279),
            .in3(N__1516),
            .lcout(\uartTxInst.rClkCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2782),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_0_LC_7_9_6 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_0_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rClkCount_0_LC_7_9_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uartTxInst.rClkCount_0_LC_7_9_6  (
            .in0(N__1321),
            .in1(N__1656),
            .in2(_gnd_net_),
            .in3(N__1518),
            .lcout(\uartTxInst.rClkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2782),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxState_RNINSDP_0_LC_7_10_0 .C_ON=1'b0;
    defparam \uartTxInst.rTxState_RNINSDP_0_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rTxState_RNINSDP_0_LC_7_10_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uartTxInst.rTxState_RNINSDP_0_LC_7_10_0  (
            .in0(N__1820),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1739),
            .lcout(\uartTxInst.rbitindex15 ),
            .ltout(\uartTxInst.rbitindex15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_1_LC_7_10_1 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_1_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rClkCount_1_LC_7_10_1 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \uartTxInst.rClkCount_1_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__1317),
            .in2(N__1402),
            .in3(N__1396),
            .lcout(\uartTxInst.rClkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2784),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_RNI85A6_5_LC_7_10_3 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_RNI85A6_5_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rClkCount_RNI85A6_5_LC_7_10_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uartTxInst.rClkCount_RNI85A6_5_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(N__1395),
            .in2(_gnd_net_),
            .in3(N__1555),
            .lcout(\uartTxInst.un2_rclkcount_5_0 ),
            .ltout(\uartTxInst.un2_rclkcount_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_RNI85BP_2_LC_7_10_4 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_RNI85BP_2_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rClkCount_RNI85BP_2_LC_7_10_4 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \uartTxInst.rClkCount_RNI85BP_2_LC_7_10_4  (
            .in0(N__1316),
            .in1(N__1740),
            .in2(N__1378),
            .in3(N__1339),
            .lcout(\uartTxInst.rTxState_10_0_x2_0_o2_d_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxDV_LC_7_10_5.C_ON=1'b0;
    defparam rTxDV_LC_7_10_5.SEQ_MODE=4'b1000;
    defparam rTxDV_LC_7_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 rTxDV_LC_7_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2300),
            .lcout(rTxDVZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2784),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_RNIOIKC_7_LC_7_10_6 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_RNIOIKC_7_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rClkCount_RNIOIKC_7_LC_7_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uartTxInst.rClkCount_RNIOIKC_7_LC_7_10_6  (
            .in0(N__1374),
            .in1(N__1577),
            .in2(N__1471),
            .in3(N__1361),
            .lcout(\uartTxInst.un2_rclkcount_4 ),
            .ltout(\uartTxInst.un2_rclkcount_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_RNI4P8P_2_LC_7_10_7 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_RNI4P8P_2_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rClkCount_RNI4P8P_2_LC_7_10_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uartTxInst.rClkCount_RNI4P8P_2_LC_7_10_7  (
            .in0(N__1338),
            .in1(N__1315),
            .in2(N__1294),
            .in3(N__1291),
            .lcout(\uartTxInst.SUM_N_3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxState_1_LC_7_11_0 .C_ON=1'b0;
    defparam \uartTxInst.rTxState_1_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rTxState_1_LC_7_11_0 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \uartTxInst.rTxState_1_LC_7_11_0  (
            .in0(N__1818),
            .in1(_gnd_net_),
            .in2(N__1755),
            .in3(N__1515),
            .lcout(\uartTxInst.rTxStateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2786),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rBitIndex_RNO_1_1_LC_7_11_1 .C_ON=1'b0;
    defparam \uartTxInst.rBitIndex_RNO_1_1_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rBitIndex_RNO_1_1_LC_7_11_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \uartTxInst.rBitIndex_RNO_1_1_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__1816),
            .in2(_gnd_net_),
            .in3(N__1901),
            .lcout(),
            .ltout(\uartTxInst.g2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rBitIndex_RNO_0_1_LC_7_11_2 .C_ON=1'b0;
    defparam \uartTxInst.rBitIndex_RNO_0_1_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rBitIndex_RNO_0_1_LC_7_11_2 .LUT_INIT=16'b0000000011110010;
    LogicCell40 \uartTxInst.rBitIndex_RNO_0_1_LC_7_11_2  (
            .in0(N__1742),
            .in1(N__1513),
            .in2(N__1441),
            .in3(N__1950),
            .lcout(),
            .ltout(\uartTxInst.rBitIndex_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rBitIndex_1_LC_7_11_3 .C_ON=1'b0;
    defparam \uartTxInst.rBitIndex_1_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rBitIndex_1_LC_7_11_3 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \uartTxInst.rBitIndex_1_LC_7_11_3  (
            .in0(N__1690),
            .in1(N__1672),
            .in2(N__1438),
            .in3(N__1699),
            .lcout(\uartTxInst.rBitIndexZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2786),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxState_RNO_1_0_LC_7_11_5 .C_ON=1'b0;
    defparam \uartTxInst.rTxState_RNO_1_0_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rTxState_RNO_1_0_LC_7_11_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uartTxInst.rTxState_RNO_1_0_LC_7_11_5  (
            .in0(N__1609),
            .in1(N__1741),
            .in2(_gnd_net_),
            .in3(N__1817),
            .lcout(\uartTxInst.rTxByte_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxState_RNO_0_0_LC_7_11_6 .C_ON=1'b0;
    defparam \uartTxInst.rTxState_RNO_0_0_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rTxState_RNO_0_0_LC_7_11_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uartTxInst.rTxState_RNO_0_0_LC_7_11_6  (
            .in0(N__1762),
            .in1(N__1842),
            .in2(N__1754),
            .in3(N__1951),
            .lcout(),
            .ltout(\uartTxInst.rTxState_10_0_i_a2_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxState_0_LC_7_11_7 .C_ON=1'b0;
    defparam \uartTxInst.rTxState_0_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rTxState_0_LC_7_11_7 .LUT_INIT=16'b1111110111101100;
    LogicCell40 \uartTxInst.rTxState_0_LC_7_11_7  (
            .in0(N__1514),
            .in1(N__1435),
            .in2(N__1429),
            .in3(N__1819),
            .lcout(\uartTxInst.rTxStateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2786),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.oSerial_LC_7_12_0 .C_ON=1'b0;
    defparam \uartTxInst.oSerial_LC_7_12_0 .SEQ_MODE=4'b1001;
    defparam \uartTxInst.oSerial_LC_7_12_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \uartTxInst.oSerial_LC_7_12_0  (
            .in0(N__1521),
            .in1(N__1750),
            .in2(N__1419),
            .in3(N__1783),
            .lcout(o_UART_TX_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2791),
            .ce(),
            .sr(N__1678));
    defparam \uartTxInst.rBitIndex_0_LC_7_12_1 .C_ON=1'b0;
    defparam \uartTxInst.rBitIndex_0_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rBitIndex_0_LC_7_12_1 .LUT_INIT=16'b1011101001000101;
    LogicCell40 \uartTxInst.rBitIndex_0_LC_7_12_1  (
            .in0(N__1822),
            .in1(N__1522),
            .in2(N__1756),
            .in3(N__1902),
            .lcout(\uartTxInst.rBitIndexZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2791),
            .ce(),
            .sr(N__1678));
    defparam CONSTANT_ONE_LUT4_LC_8_8_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_8_8_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_8_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_RNO_0_6_LC_8_9_1 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_RNO_0_6_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rClkCount_RNO_0_6_LC_8_9_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uartTxInst.rClkCount_RNO_0_6_LC_8_9_1  (
            .in0(N__1578),
            .in1(N__1556),
            .in2(N__1537),
            .in3(N__1464),
            .lcout(),
            .ltout(\uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_6_LC_8_9_2 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_6_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rClkCount_6_LC_8_9_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \uartTxInst.rClkCount_6_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__1517),
            .in2(N__1582),
            .in3(N__1666),
            .lcout(\uartTxInst.rClkCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2785),
            .ce(),
            .sr(_gnd_net_));
    defparam rRamAddress_0_LC_8_9_3.C_ON=1'b0;
    defparam rRamAddress_0_LC_8_9_3.SEQ_MODE=4'b1000;
    defparam rRamAddress_0_LC_8_9_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 rRamAddress_0_LC_8_9_3 (
            .in0(N__2299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2253),
            .lcout(rRamAddressZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2785),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_5_LC_8_9_4 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_5_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rClkCount_5_LC_8_9_4 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \uartTxInst.rClkCount_5_LC_8_9_4  (
            .in0(N__1465),
            .in1(N__1665),
            .in2(N__1561),
            .in3(N__1536),
            .lcout(\uartTxInst.rClkCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2785),
            .ce(),
            .sr(_gnd_net_));
    defparam rRamAddress_2_LC_8_9_5.C_ON=1'b0;
    defparam rRamAddress_2_LC_8_9_5.SEQ_MODE=4'b1000;
    defparam rRamAddress_2_LC_8_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRamAddress_2_LC_8_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2169),
            .lcout(rRamAddressZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2785),
            .ce(),
            .sr(_gnd_net_));
    defparam rRamAddress_1_LC_8_9_6.C_ON=1'b0;
    defparam rRamAddress_1_LC_8_9_6.SEQ_MODE=4'b1000;
    defparam rRamAddress_1_LC_8_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRamAddress_1_LC_8_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2205),
            .lcout(rRamAddressZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2785),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rClkCount_4_LC_8_9_7 .C_ON=1'b0;
    defparam \uartTxInst.rClkCount_4_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rClkCount_4_LC_8_9_7 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \uartTxInst.rClkCount_4_LC_8_9_7  (
            .in0(N__1535),
            .in1(N__1466),
            .in2(N__1677),
            .in3(N__1520),
            .lcout(\uartTxInst.rClkCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2785),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxByte_7_LC_8_10_0 .C_ON=1'b0;
    defparam \uartTxInst.rTxByte_7_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rTxByte_7_LC_8_10_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \uartTxInst.rTxByte_7_LC_8_10_0  (
            .in0(N__1671),
            .in1(N__1608),
            .in2(N__2317),
            .in3(N__1873),
            .lcout(\uartTxInst.rTxByte_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2787),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxByte_4_LC_8_10_1 .C_ON=1'b0;
    defparam \uartTxInst.rTxByte_4_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rTxByte_4_LC_8_10_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \uartTxInst.rTxByte_4_LC_8_10_1  (
            .in0(N__1605),
            .in1(N__1668),
            .in2(N__2365),
            .in3(N__1929),
            .lcout(\uartTxInst.rTxByte_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2787),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxByte_6_LC_8_10_2 .C_ON=1'b0;
    defparam \uartTxInst.rTxByte_6_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rTxByte_6_LC_8_10_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \uartTxInst.rTxByte_6_LC_8_10_2  (
            .in0(N__1670),
            .in1(N__1607),
            .in2(N__2335),
            .in3(N__1915),
            .lcout(\uartTxInst.rTxByte_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2787),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rBitIndex_RNI0NON_0_LC_8_10_3 .C_ON=1'b0;
    defparam \uartTxInst.rBitIndex_RNI0NON_0_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rBitIndex_RNI0NON_0_LC_8_10_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \uartTxInst.rBitIndex_RNI0NON_0_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__1815),
            .in2(_gnd_net_),
            .in3(N__1903),
            .lcout(\uartTxInst.N_31 ),
            .ltout(\uartTxInst.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rBitIndex_RNIQ26S1_1_LC_8_10_4 .C_ON=1'b0;
    defparam \uartTxInst.rBitIndex_RNIQ26S1_1_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.rBitIndex_RNIQ26S1_1_LC_8_10_4 .LUT_INIT=16'b1111001011111111;
    LogicCell40 \uartTxInst.rBitIndex_RNIQ26S1_1_LC_8_10_4  (
            .in0(N__1749),
            .in1(N__1708),
            .in2(N__1702),
            .in3(N__1949),
            .lcout(\uartTxInst.rTxState_10_0_x2_0_o2_1_1_1 ),
            .ltout(\uartTxInst.rTxState_10_0_x2_0_o2_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rBitIndex_2_LC_8_10_5 .C_ON=1'b0;
    defparam \uartTxInst.rBitIndex_2_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rBitIndex_2_LC_8_10_5 .LUT_INIT=16'b0010001000100001;
    LogicCell40 \uartTxInst.rBitIndex_2_LC_8_10_5  (
            .in0(N__1843),
            .in1(N__1667),
            .in2(N__1693),
            .in3(N__1689),
            .lcout(\uartTxInst.rBitIndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2787),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.rTxByte_5_LC_8_10_6 .C_ON=1'b0;
    defparam \uartTxInst.rTxByte_5_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \uartTxInst.rTxByte_5_LC_8_10_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \uartTxInst.rTxByte_5_LC_8_10_6  (
            .in0(N__1669),
            .in1(N__1606),
            .in2(N__1858),
            .in3(N__2347),
            .lcout(\uartTxInst.rTxByte_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2787),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rDataReady_LC_8_10_7 .C_ON=1'b0;
    defparam \uartRxInst.rDataReady_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rDataReady_LC_8_10_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \uartRxInst.rDataReady_LC_8_10_7  (
            .in0(N__2916),
            .in1(N__3047),
            .in2(_gnd_net_),
            .in3(N__2298),
            .lcout(rRxReady),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2787),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rDataCounter_RNO_0_1_LC_8_11_0 .C_ON=1'b0;
    defparam \uartRxInst.rDataCounter_RNO_0_1_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rDataCounter_RNO_0_1_LC_8_11_0 .LUT_INIT=16'b1101001011110000;
    LogicCell40 \uartRxInst.rDataCounter_RNO_0_1_LC_8_11_0  (
            .in0(N__2081),
            .in1(N__3043),
            .in2(N__2104),
            .in3(N__2491),
            .lcout(),
            .ltout(\uartRxInst.rDataCounter_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rDataCounter_1_LC_8_11_1 .C_ON=1'b0;
    defparam \uartRxInst.rDataCounter_1_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rDataCounter_1_LC_8_11_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uartRxInst.rDataCounter_1_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1585),
            .in3(N__2459),
            .lcout(\uartRxInst.rDataCounterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2792),
            .ce(),
            .sr(N__2443));
    defparam \uartRxInst.rDataCounter_0_LC_8_11_2 .C_ON=1'b0;
    defparam \uartRxInst.rDataCounter_0_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rDataCounter_0_LC_8_11_2 .LUT_INIT=16'b1111100111111010;
    LogicCell40 \uartRxInst.rDataCounter_0_LC_8_11_2  (
            .in0(N__2082),
            .in1(N__3044),
            .in2(N__2464),
            .in3(N__2492),
            .lcout(\uartRxInst.rDataCounterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2792),
            .ce(),
            .sr(N__2443));
    defparam \uartRxInst.rDataCounter_RNILM1D1_2_LC_8_11_3 .C_ON=1'b0;
    defparam \uartRxInst.rDataCounter_RNILM1D1_2_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rDataCounter_RNILM1D1_2_LC_8_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uartRxInst.rDataCounter_RNILM1D1_2_LC_8_11_3  (
            .in0(N__1773),
            .in1(N__2099),
            .in2(_gnd_net_),
            .in3(N__2080),
            .lcout(\uartRxInst.rState_0_sqmuxa_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.oSerial_RNO_2_LC_8_11_4 .C_ON=1'b0;
    defparam \uartTxInst.oSerial_RNO_2_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.oSerial_RNO_2_LC_8_11_4 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \uartTxInst.oSerial_RNO_2_LC_8_11_4  (
            .in0(N__1948),
            .in1(N__1899),
            .in2(N__1930),
            .in3(N__1914),
            .lcout(),
            .ltout(\uartTxInst.oSerial_3_6_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.oSerial_RNO_1_LC_8_11_5 .C_ON=1'b0;
    defparam \uartTxInst.oSerial_RNO_1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.oSerial_RNO_1_LC_8_11_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \uartTxInst.oSerial_RNO_1_LC_8_11_5  (
            .in0(N__1900),
            .in1(N__1872),
            .in2(N__1861),
            .in3(N__1854),
            .lcout(),
            .ltout(\uartTxInst.N_35_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartTxInst.oSerial_RNO_0_LC_8_11_6 .C_ON=1'b0;
    defparam \uartTxInst.oSerial_RNO_0_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \uartTxInst.oSerial_RNO_0_LC_8_11_6 .LUT_INIT=16'b0000000000111111;
    LogicCell40 \uartTxInst.oSerial_RNO_0_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__1841),
            .in2(N__1825),
            .in3(N__1821),
            .lcout(\uartTxInst.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rDataCounter_2_LC_8_11_7 .C_ON=1'b0;
    defparam \uartRxInst.rDataCounter_2_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rDataCounter_2_LC_8_11_7 .LUT_INIT=16'b1111111101111000;
    LogicCell40 \uartRxInst.rDataCounter_2_LC_8_11_7  (
            .in0(N__2493),
            .in1(N__2065),
            .in2(N__1777),
            .in3(N__2463),
            .lcout(\uartRxInst.rDataCounterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2792),
            .ce(),
            .sr(N__2443));
    defparam \uartRxInst.rCycleCounter_RNI66KJ1_7_LC_8_12_0 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_RNI66KJ1_7_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNI66KJ1_7_LC_8_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uartRxInst.rCycleCounter_RNI66KJ1_7_LC_8_12_0  (
            .in0(N__2517),
            .in1(N__2684),
            .in2(N__2548),
            .in3(N__2633),
            .lcout(\uartRxInst.g0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rState_RNIRJB_0_1_LC_8_12_1 .C_ON=1'b0;
    defparam \uartRxInst.rState_RNIRJB_0_1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rState_RNIRJB_0_1_LC_8_12_1 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uartRxInst.rState_RNIRJB_0_1_LC_8_12_1  (
            .in0(N__3041),
            .in1(N__2910),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uartRxInst.rstateZ0 ),
            .ltout(\uartRxInst.rstateZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_5_LC_8_12_2 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_5_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rCycleCounter_5_LC_8_12_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \uartRxInst.rCycleCounter_5_LC_8_12_2  (
            .in0(N__2979),
            .in1(N__2848),
            .in2(N__1765),
            .in3(N__2041),
            .lcout(\uartRxInst.rCycleCounterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2794),
            .ce(N__2735),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_6_LC_8_12_3 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_6_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rCycleCounter_6_LC_8_12_3 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \uartRxInst.rCycleCounter_6_LC_8_12_3  (
            .in0(N__2849),
            .in1(N__2980),
            .in2(N__2926),
            .in3(N__1960),
            .lcout(\uartRxInst.rCycleCounterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2794),
            .ce(N__2735),
            .sr(_gnd_net_));
    defparam \uartRxInst.rState_RNIRJB_1_LC_8_12_5 .C_ON=1'b0;
    defparam \uartRxInst.rState_RNIRJB_1_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rState_RNIRJB_1_LC_8_12_5 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \uartRxInst.rState_RNIRJB_1_LC_8_12_5  (
            .in0(N__3042),
            .in1(N__2909),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uartRxInst.rCycleCountere_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_4_LC_8_12_6 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_4_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rCycleCounter_4_LC_8_12_6 .LUT_INIT=16'b0010111000011101;
    LogicCell40 \uartRxInst.rCycleCounter_4_LC_8_12_6  (
            .in0(N__2518),
            .in1(N__2850),
            .in2(N__2584),
            .in3(N__2050),
            .lcout(\uartRxInst.rCycleCounterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2794),
            .ce(N__2735),
            .sr(_gnd_net_));
    defparam \uartRxInst.rDataCounter_RNO_0_2_LC_8_12_7 .C_ON=1'b0;
    defparam \uartRxInst.rDataCounter_RNO_0_2_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rDataCounter_RNO_0_2_LC_8_12_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uartRxInst.rDataCounter_RNO_0_2_LC_8_12_7  (
            .in0(N__3040),
            .in1(N__2103),
            .in2(_gnd_net_),
            .in3(N__2086),
            .lcout(\uartRxInst.CO1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_cry_c_0_LC_8_13_0 .C_ON=1'b1;
    defparam \uartRxInst.rCycleCounter_cry_c_0_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_cry_c_0_LC_8_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uartRxInst.rCycleCounter_cry_c_0_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__2820),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\uartRxInst.rCycleCounter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_cry_0_THRU_LUT4_0_LC_8_13_1 .C_ON=1'b1;
    defparam \uartRxInst.rCycleCounter_cry_0_THRU_LUT4_0_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_cry_0_THRU_LUT4_0_LC_8_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uartRxInst.rCycleCounter_cry_0_THRU_LUT4_0_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__3077),
            .in2(N__2020),
            .in3(N__2059),
            .lcout(\uartRxInst.rCycleCounter_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\uartRxInst.rCycleCounter_cry_0 ),
            .carryout(\uartRxInst.rCycleCounter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNO_0_2_LC_8_13_2 .C_ON=1'b1;
    defparam \uartRxInst.rCycleCounter_RNO_0_2_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNO_0_2_LC_8_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uartRxInst.rCycleCounter_RNO_0_2_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__2709),
            .in2(N__2030),
            .in3(N__2056),
            .lcout(\uartRxInst.rCycleCounter_s_2 ),
            .ltout(),
            .carryin(\uartRxInst.rCycleCounter_cry_1 ),
            .carryout(\uartRxInst.rCycleCounter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNO_0_3_LC_8_13_3 .C_ON=1'b1;
    defparam \uartRxInst.rCycleCounter_RNO_0_3_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNO_0_3_LC_8_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uartRxInst.rCycleCounter_RNO_0_3_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__2660),
            .in2(N__2018),
            .in3(N__2053),
            .lcout(\uartRxInst.rCycleCounter_s_3 ),
            .ltout(),
            .carryin(\uartRxInst.rCycleCounter_cry_2 ),
            .carryout(\uartRxInst.rCycleCounter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_cry_3_THRU_LUT4_0_LC_8_13_4 .C_ON=1'b1;
    defparam \uartRxInst.rCycleCounter_cry_3_THRU_LUT4_0_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_cry_3_THRU_LUT4_0_LC_8_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uartRxInst.rCycleCounter_cry_3_THRU_LUT4_0_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__2521),
            .in2(N__2032),
            .in3(N__2044),
            .lcout(\uartRxInst.rCycleCounter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\uartRxInst.rCycleCounter_cry_3 ),
            .carryout(\uartRxInst.rCycleCounter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNO_0_5_LC_8_13_5 .C_ON=1'b1;
    defparam \uartRxInst.rCycleCounter_RNO_0_5_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNO_0_5_LC_8_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uartRxInst.rCycleCounter_RNO_0_5_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__2547),
            .in2(N__2019),
            .in3(N__2035),
            .lcout(\uartRxInst.rCycleCounter_s_5 ),
            .ltout(),
            .carryin(\uartRxInst.rCycleCounter_cry_4 ),
            .carryout(\uartRxInst.rCycleCounter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNO_0_6_LC_8_13_6 .C_ON=1'b1;
    defparam \uartRxInst.rCycleCounter_RNO_0_6_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNO_0_6_LC_8_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uartRxInst.rCycleCounter_RNO_0_6_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__2635),
            .in2(N__2031),
            .in3(N__1954),
            .lcout(\uartRxInst.rCycleCounter_s_6 ),
            .ltout(),
            .carryin(\uartRxInst.rCycleCounter_cry_5 ),
            .carryout(\uartRxInst.rCycleCounter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_7_LC_8_13_7 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_7_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rCycleCounter_7_LC_8_13_7 .LUT_INIT=16'b0111010001000111;
    LogicCell40 \uartRxInst.rCycleCounter_7_LC_8_13_7  (
            .in0(N__2580),
            .in1(N__2851),
            .in2(N__2689),
            .in3(N__2263),
            .lcout(\uartRxInst.rCycleCounterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2796),
            .ce(N__2742),
            .sr(_gnd_net_));
    defparam rRamAddress_4_LC_9_8_6.C_ON=1'b0;
    defparam rRamAddress_4_LC_9_8_6.SEQ_MODE=4'b1000;
    defparam rRamAddress_4_LC_9_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRamAddress_4_LC_9_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2130),
            .lcout(rRamAddressZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2783),
            .ce(),
            .sr(_gnd_net_));
    defparam rRamAddress_RNIJ99L_0_LC_9_9_0.C_ON=1'b1;
    defparam rRamAddress_RNIJ99L_0_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam rRamAddress_RNIJ99L_0_LC_9_9_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 rRamAddress_RNIJ99L_0_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(N__2252),
            .in2(N__2304),
            .in3(N__2297),
            .lcout(pEcho_rRamAddress_2_0),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(pEcho_rRamAddress_2_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pEcho_rRamAddress_2_cry_0_c_RNI5QRQ_LC_9_9_1.C_ON=1'b1;
    defparam pEcho_rRamAddress_2_cry_0_c_RNI5QRQ_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam pEcho_rRamAddress_2_cry_0_c_RNI5QRQ_LC_9_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 pEcho_rRamAddress_2_cry_0_c_RNI5QRQ_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(N__2220),
            .in2(_gnd_net_),
            .in3(N__2194),
            .lcout(pEcho_rRamAddress_2_1),
            .ltout(),
            .carryin(pEcho_rRamAddress_2_cry_0),
            .carryout(pEcho_rRamAddress_2_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pEcho_rRamAddress_2_cry_1_c_RNI7TSQ_LC_9_9_2.C_ON=1'b1;
    defparam pEcho_rRamAddress_2_cry_1_c_RNI7TSQ_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam pEcho_rRamAddress_2_cry_1_c_RNI7TSQ_LC_9_9_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 pEcho_rRamAddress_2_cry_1_c_RNI7TSQ_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(N__2184),
            .in2(_gnd_net_),
            .in3(N__2158),
            .lcout(pEcho_rRamAddress_2_2),
            .ltout(),
            .carryin(pEcho_rRamAddress_2_cry_1),
            .carryout(pEcho_rRamAddress_2_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pEcho_rRamAddress_2_cry_2_c_RNI90UQ_LC_9_9_3.C_ON=1'b1;
    defparam pEcho_rRamAddress_2_cry_2_c_RNI90UQ_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam pEcho_rRamAddress_2_cry_2_c_RNI90UQ_LC_9_9_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 pEcho_rRamAddress_2_cry_2_c_RNI90UQ_LC_9_9_3 (
            .in0(_gnd_net_),
            .in1(N__2382),
            .in2(_gnd_net_),
            .in3(N__2155),
            .lcout(pEcho_rRamAddress_2_3),
            .ltout(),
            .carryin(pEcho_rRamAddress_2_cry_2),
            .carryout(pEcho_rRamAddress_2_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pEcho_rRamAddress_2_cry_3_c_RNIB3VQ_LC_9_9_4.C_ON=1'b1;
    defparam pEcho_rRamAddress_2_cry_3_c_RNIB3VQ_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam pEcho_rRamAddress_2_cry_3_c_RNIB3VQ_LC_9_9_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 pEcho_rRamAddress_2_cry_3_c_RNIB3VQ_LC_9_9_4 (
            .in0(_gnd_net_),
            .in1(N__2145),
            .in2(_gnd_net_),
            .in3(N__2119),
            .lcout(pEcho_rRamAddress_2_4),
            .ltout(),
            .carryin(pEcho_rRamAddress_2_cry_3),
            .carryout(pEcho_rRamAddress_2_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pEcho_rRamAddress_2_cry_4_c_RNID60R_LC_9_9_5.C_ON=1'b0;
    defparam pEcho_rRamAddress_2_cry_4_c_RNID60R_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam pEcho_rRamAddress_2_cry_4_c_RNID60R_LC_9_9_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 pEcho_rRamAddress_2_cry_4_c_RNID60R_LC_9_9_5 (
            .in0(_gnd_net_),
            .in1(N__2412),
            .in2(_gnd_net_),
            .in3(N__2116),
            .lcout(pEcho_rRamAddress_2_5),
            .ltout(pEcho_rRamAddress_2_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rRamAddress_5_LC_9_9_6.C_ON=1'b0;
    defparam rRamAddress_5_LC_9_9_6.SEQ_MODE=4'b1000;
    defparam rRamAddress_5_LC_9_9_6.LUT_INIT=16'b1111000011110000;
    LogicCell40 rRamAddress_5_LC_9_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2419),
            .in3(_gnd_net_),
            .lcout(rRamAddressZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2788),
            .ce(),
            .sr(_gnd_net_));
    defparam rRamAddress_3_LC_9_9_7.C_ON=1'b0;
    defparam rRamAddress_3_LC_9_9_7.SEQ_MODE=4'b1000;
    defparam rRamAddress_3_LC_9_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRamAddress_3_LC_9_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2397),
            .lcout(rRamAddressZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2788),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_e_0_4_LC_9_10_0.C_ON=1'b0;
    defparam rTxByte_e_0_4_LC_9_10_0.SEQ_MODE=4'b1000;
    defparam rTxByte_e_0_4_LC_9_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 rTxByte_e_0_4_LC_9_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2371),
            .lcout(rTxByteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2793),
            .ce(N__2305),
            .sr(_gnd_net_));
    defparam rTxByte_e_0_5_LC_9_10_1.C_ON=1'b0;
    defparam rTxByte_e_0_5_LC_9_10_1.SEQ_MODE=4'b1000;
    defparam rTxByte_e_0_5_LC_9_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 rTxByte_e_0_5_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2353),
            .lcout(rTxByteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2793),
            .ce(N__2305),
            .sr(_gnd_net_));
    defparam rTxByte_e_0_6_LC_9_10_2.C_ON=1'b0;
    defparam rTxByte_e_0_6_LC_9_10_2.SEQ_MODE=4'b1000;
    defparam rTxByte_e_0_6_LC_9_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 rTxByte_e_0_6_LC_9_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2341),
            .lcout(rTxByteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2793),
            .ce(N__2305),
            .sr(_gnd_net_));
    defparam rTxByte_e_0_7_LC_9_10_3.C_ON=1'b0;
    defparam rTxByte_e_0_7_LC_9_10_3.SEQ_MODE=4'b1000;
    defparam rTxByte_e_0_7_LC_9_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 rTxByte_e_0_7_LC_9_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2323),
            .lcout(rTxByteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2793),
            .ce(N__2305),
            .sr(_gnd_net_));
    defparam \uartRxInst.rState_1_LC_9_11_0 .C_ON=1'b0;
    defparam \uartRxInst.rState_1_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rState_1_LC_9_11_0 .LUT_INIT=16'b0001000111001100;
    LogicCell40 \uartRxInst.rState_1_LC_9_11_0  (
            .in0(N__2983),
            .in1(N__2918),
            .in2(_gnd_net_),
            .in3(N__3046),
            .lcout(uartRxInst_rState_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2795),
            .ce(N__2560),
            .sr(_gnd_net_));
    defparam \uartRxInst.rState_0_LC_9_11_2 .C_ON=1'b0;
    defparam \uartRxInst.rState_0_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rState_0_LC_9_11_2 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uartRxInst.rState_0_LC_9_11_2  (
            .in0(N__2982),
            .in1(N__2917),
            .in2(_gnd_net_),
            .in3(N__3045),
            .lcout(uartRxInst_rState_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2795),
            .ce(N__2560),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNICOS61_1_LC_9_12_0 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_RNICOS61_1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNICOS61_1_LC_9_12_0 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \uartRxInst.rCycleCounter_RNICOS61_1_LC_9_12_0  (
            .in0(N__2545),
            .in1(N__2520),
            .in2(N__2922),
            .in3(N__3076),
            .lcout(G_11_i_a3_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNIAMVP_0_LC_9_12_1 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_RNIAMVP_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNIAMVP_0_LC_9_12_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uartRxInst.rCycleCounter_RNIAMVP_0_LC_9_12_1  (
            .in0(N__3048),
            .in1(N__2544),
            .in2(_gnd_net_),
            .in3(N__2821),
            .lcout(),
            .ltout(G_11_i_a3_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i_UART_RX_ibuf_RNI5MUN3_LC_9_12_2.C_ON=1'b0;
    defparam i_UART_RX_ibuf_RNI5MUN3_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam i_UART_RX_ibuf_RNI5MUN3_LC_9_12_2.LUT_INIT=16'b0001010101010101;
    LogicCell40 i_UART_RX_ibuf_RNI5MUN3_LC_9_12_2 (
            .in0(N__2569),
            .in1(N__2593),
            .in2(N__2587),
            .in3(N__2611),
            .lcout(uartRxInst_un1_rData_0_sqmuxa_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i_UART_RX_ibuf_RNID5E3_LC_9_12_3.C_ON=1'b0;
    defparam i_UART_RX_ibuf_RNID5E3_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam i_UART_RX_ibuf_RNID5E3_LC_9_12_3.LUT_INIT=16'b0000000000100010;
    LogicCell40 i_UART_RX_ibuf_RNID5E3_LC_9_12_3 (
            .in0(N__3049),
            .in1(N__2901),
            .in2(_gnd_net_),
            .in3(N__2978),
            .lcout(N_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rState_RNIC6LK4_1_LC_9_12_4 .C_ON=1'b0;
    defparam \uartRxInst.rState_RNIC6LK4_1_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rState_RNIC6LK4_1_LC_9_12_4 .LUT_INIT=16'b1110111111000011;
    LogicCell40 \uartRxInst.rState_RNIC6LK4_1_LC_9_12_4  (
            .in0(N__2473),
            .in1(N__3051),
            .in2(N__2923),
            .in3(N__2494),
            .lcout(\uartRxInst.un1_rCycleCounter_2_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNI55QP_7_LC_9_12_5 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_RNI55QP_7_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNI55QP_7_LC_9_12_5 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \uartRxInst.rCycleCounter_RNI55QP_7_LC_9_12_5  (
            .in0(N__2683),
            .in1(N__2632),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\uartRxInst.un12_rstate_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNISR773_4_LC_9_12_6 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_RNISR773_4_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNISR773_4_LC_9_12_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uartRxInst.rCycleCounter_RNISR773_4_LC_9_12_6  (
            .in0(N__2546),
            .in1(N__2519),
            .in2(N__2497),
            .in3(N__3088),
            .lcout(\uartRxInst.N_83_0_i ),
            .ltout(\uartRxInst.N_83_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rState_RNIC6LK4_0_1_LC_9_12_7 .C_ON=1'b0;
    defparam \uartRxInst.rState_RNIC6LK4_0_1_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rState_RNIC6LK4_0_1_LC_9_12_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uartRxInst.rState_RNIC6LK4_0_1_LC_9_12_7  (
            .in0(N__3050),
            .in1(N__2908),
            .in2(N__2476),
            .in3(N__2472),
            .lcout(\uartRxInst.rDataCounter_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_1_LC_9_13_0 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_1_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rCycleCounter_1_LC_9_13_0 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \uartRxInst.rCycleCounter_1_LC_9_13_0  (
            .in0(N__2847),
            .in1(N__2449),
            .in2(_gnd_net_),
            .in3(N__3081),
            .lcout(\uartRxInst.rCycleCounterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2797),
            .ce(N__2743),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_2_LC_9_13_1 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_2_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rCycleCounter_2_LC_9_13_1 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \uartRxInst.rCycleCounter_2_LC_9_13_1  (
            .in0(N__2442),
            .in1(N__2425),
            .in2(N__2981),
            .in3(N__2845),
            .lcout(\uartRxInst.rCycleCounterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2797),
            .ce(N__2743),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNIMLJJ1_0_0_LC_9_13_2 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_RNIMLJJ1_0_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNIMLJJ1_0_0_LC_9_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uartRxInst.rCycleCounter_RNIMLJJ1_0_0_LC_9_13_2  (
            .in0(N__3075),
            .in1(N__2817),
            .in2(N__2661),
            .in3(N__2707),
            .lcout(\uartRxInst.un12_rstate_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNIMLJJ1_0_LC_9_13_3 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_RNIMLJJ1_0_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNIMLJJ1_0_LC_9_13_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uartRxInst.rCycleCounter_RNIMLJJ1_0_LC_9_13_3  (
            .in0(N__2818),
            .in1(N__2656),
            .in2(N__3082),
            .in3(N__2710),
            .lcout(),
            .ltout(\uartRxInst.g0_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rState_RNINFJ73_1_LC_9_13_4 .C_ON=1'b0;
    defparam \uartRxInst.rState_RNINFJ73_1_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rState_RNINFJ73_1_LC_9_13_4 .LUT_INIT=16'b1111000100010001;
    LogicCell40 \uartRxInst.rState_RNINFJ73_1_LC_9_13_4  (
            .in0(N__2924),
            .in1(N__3052),
            .in2(N__2992),
            .in3(N__2989),
            .lcout(\uartRxInst.N_83_0_i_0 ),
            .ltout(\uartRxInst.N_83_0_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_3_LC_9_13_5 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_3_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rCycleCounter_3_LC_9_13_5 .LUT_INIT=16'b1101111111010000;
    LogicCell40 \uartRxInst.rCycleCounter_3_LC_9_13_5  (
            .in0(N__2972),
            .in1(N__2925),
            .in2(N__2860),
            .in3(N__2857),
            .lcout(\uartRxInst.rCycleCounterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2797),
            .ce(N__2743),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_0_LC_9_13_6 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_0_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \uartRxInst.rCycleCounter_0_LC_9_13_6 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \uartRxInst.rCycleCounter_0_LC_9_13_6  (
            .in0(N__2846),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2819),
            .lcout(\uartRxInst.rCycleCounterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2797),
            .ce(N__2743),
            .sr(_gnd_net_));
    defparam \uartRxInst.rCycleCounter_RNI22KJ1_7_LC_9_13_7 .C_ON=1'b0;
    defparam \uartRxInst.rCycleCounter_RNI22KJ1_7_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \uartRxInst.rCycleCounter_RNI22KJ1_7_LC_9_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uartRxInst.rCycleCounter_RNI22KJ1_7_LC_9_13_7  (
            .in0(N__2708),
            .in1(N__2685),
            .in2(N__2662),
            .in3(N__2634),
            .lcout(G_11_i_a3_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ZERO_LUT4_LC_11_9_0.C_ON=1'b0;
    defparam CONSTANT_ZERO_LUT4_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ZERO_LUT4_LC_11_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 CONSTANT_ZERO_LUT4_LC_11_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ZERO_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // core
