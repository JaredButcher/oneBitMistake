-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 28 2019 14:20:42

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "core" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of core
entity core is
port (
    o_UART_TX : out std_logic;
    i_UART_RX : in std_logic;
    i_Clk : in std_logic);
end core;

-- Architecture of core
-- View name is \INTERFACE\
architecture \INTERFACE\ of core is

signal \N__3127\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2170\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2124\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2082\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2062\ : std_logic;
signal \N__2059\ : std_logic;
signal \N__2056\ : std_logic;
signal \N__2053\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2047\ : std_logic;
signal \N__2044\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2032\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2019\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2011\ : std_logic;
signal \N__2010\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1997\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1984\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1973\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1951\ : std_logic;
signal \N__1950\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1930\ : std_logic;
signal \N__1929\ : std_logic;
signal \N__1926\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1920\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1914\ : std_logic;
signal \N__1911\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1902\ : std_logic;
signal \N__1901\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1899\ : std_logic;
signal \N__1896\ : std_logic;
signal \N__1893\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1866\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1854\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1841\ : std_logic;
signal \N__1838\ : std_logic;
signal \N__1835\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1821\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1818\ : std_logic;
signal \N__1817\ : std_logic;
signal \N__1816\ : std_logic;
signal \N__1815\ : std_logic;
signal \N__1812\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1806\ : std_logic;
signal \N__1797\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1783\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1777\ : std_logic;
signal \N__1774\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1755\ : std_logic;
signal \N__1754\ : std_logic;
signal \N__1751\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1746\ : std_logic;
signal \N__1743\ : std_logic;
signal \N__1742\ : std_logic;
signal \N__1741\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1739\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1722\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1708\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1690\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1683\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1677\ : std_logic;
signal \N__1676\ : std_logic;
signal \N__1673\ : std_logic;
signal \N__1672\ : std_logic;
signal \N__1671\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1666\ : std_logic;
signal \N__1665\ : std_logic;
signal \N__1662\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1660\ : std_logic;
signal \N__1657\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1650\ : std_logic;
signal \N__1639\ : std_logic;
signal \N__1632\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1622\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1608\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1590\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1574\ : std_logic;
signal \N__1571\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1560\ : std_logic;
signal \N__1557\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1537\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1525\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1521\ : std_logic;
signal \N__1520\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1518\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1515\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1494\ : std_logic;
signal \N__1487\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1468\ : std_logic;
signal \N__1467\ : std_logic;
signal \N__1466\ : std_logic;
signal \N__1465\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1461\ : std_logic;
signal \N__1458\ : std_logic;
signal \N__1451\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1441\ : std_logic;
signal \N__1438\ : std_logic;
signal \N__1435\ : std_logic;
signal \N__1432\ : std_logic;
signal \N__1429\ : std_logic;
signal \N__1426\ : std_logic;
signal \N__1423\ : std_logic;
signal \N__1420\ : std_logic;
signal \N__1419\ : std_logic;
signal \N__1416\ : std_logic;
signal \N__1413\ : std_logic;
signal \N__1410\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1402\ : std_logic;
signal \N__1399\ : std_logic;
signal \N__1398\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1396\ : std_logic;
signal \N__1395\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1383\ : std_logic;
signal \N__1378\ : std_logic;
signal \N__1375\ : std_logic;
signal \N__1374\ : std_logic;
signal \N__1371\ : std_logic;
signal \N__1368\ : std_logic;
signal \N__1363\ : std_logic;
signal \N__1362\ : std_logic;
signal \N__1361\ : std_logic;
signal \N__1356\ : std_logic;
signal \N__1353\ : std_logic;
signal \N__1348\ : std_logic;
signal \N__1347\ : std_logic;
signal \N__1346\ : std_logic;
signal \N__1343\ : std_logic;
signal \N__1340\ : std_logic;
signal \N__1339\ : std_logic;
signal \N__1338\ : std_logic;
signal \N__1331\ : std_logic;
signal \N__1326\ : std_logic;
signal \N__1321\ : std_logic;
signal \N__1320\ : std_logic;
signal \N__1319\ : std_logic;
signal \N__1318\ : std_logic;
signal \N__1317\ : std_logic;
signal \N__1316\ : std_logic;
signal \N__1315\ : std_logic;
signal \N__1306\ : std_logic;
signal \N__1299\ : std_logic;
signal \N__1294\ : std_logic;
signal \N__1291\ : std_logic;
signal \N__1288\ : std_logic;
signal \N__1285\ : std_logic;
signal \N__1282\ : std_logic;
signal \N__1279\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uartTxInst.un5_rclkcount_c4_cascade_\ : std_logic;
signal \uartTxInst.un5_rclkcount_ac0_11_cascade_\ : std_logic;
signal \uartTxInst.un5_rclkcount_c3_cascade_\ : std_logic;
signal \uartTxInst.rbitindex15_cascade_\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_1\ : std_logic;
signal \uartTxInst.un2_rclkcount_5_0_cascade_\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_7\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_3\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_2\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_0\ : std_logic;
signal \uartTxInst.un2_rclkcount_4_cascade_\ : std_logic;
signal \uartTxInst.un2_rclkcount_5_0\ : std_logic;
signal \uartTxInst.g2_0_cascade_\ : std_logic;
signal \uartTxInst.rBitIndex_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \uartTxInst.rTxByte_0_sqmuxa\ : std_logic;
signal \uartTxInst.rTxState_10_0_i_a2_1_2_0_cascade_\ : std_logic;
signal \o_UART_TX_c\ : std_logic;
signal \uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_6\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_5\ : std_logic;
signal \uartTxInst.un5_rclkcount_c4\ : std_logic;
signal \uartTxInst.SUM_N_3_mux\ : std_logic;
signal \uartTxInst.rClkCountZ0Z_4\ : std_logic;
signal \uartTxInst.N_31\ : std_logic;
signal \uartTxInst.rTxStateZ0Z_1\ : std_logic;
signal \uartTxInst.un2_rclkcount_4\ : std_logic;
signal \uartTxInst.N_31_cascade_\ : std_logic;
signal \uartTxInst.rTxState_10_0_x2_0_o2_1_1_1\ : std_logic;
signal \uartTxInst.rTxState_10_0_x2_0_o2_1_1_1_cascade_\ : std_logic;
signal \uartTxInst.rTxState_10_0_x2_0_o2_d_0_1\ : std_logic;
signal \uartTxInst.rbitindex15\ : std_logic;
signal \rTxDVZ0\ : std_logic;
signal \uartRxInst.rDataCounter_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \uartTxInst.rBitIndexZ0Z_1\ : std_logic;
signal \uartTxInst.rTxByte_0_4\ : std_logic;
signal \uartTxInst.rTxByte_0_6\ : std_logic;
signal \uartTxInst.rBitIndexZ1Z_0\ : std_logic;
signal \uartTxInst.rTxByte_0_7\ : std_logic;
signal \uartTxInst.oSerial_3_6_i_m2_ns_1_cascade_\ : std_logic;
signal \uartTxInst.rTxByte_0_5\ : std_logic;
signal \uartTxInst.rBitIndexZ0Z_2\ : std_logic;
signal \uartTxInst.N_35_cascade_\ : std_logic;
signal \uartTxInst.rTxStateZ0Z_0\ : std_logic;
signal \uartTxInst.N_48\ : std_logic;
signal \uartRxInst.rDataCounterZ0Z_2\ : std_logic;
signal \uartRxInst.rstateZ0_cascade_\ : std_logic;
signal \uartRxInst.rDataCounterZ0Z_1\ : std_logic;
signal \uartRxInst.rDataCounterZ0Z_0\ : std_logic;
signal \uartRxInst.CO1_0\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_0\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_1\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_2\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_3_THRU_CO\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_3\ : std_logic;
signal \uartRxInst.rCycleCounter_s_5\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_4\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \uartRxInst.rCycleCounter_s_6\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_5\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_6\ : std_logic;
signal \rRamAddressZ0Z_0\ : std_logic;
signal \pEcho_rRamAddress_2_0\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \rRamAddressZ0Z_1\ : std_logic;
signal \pEcho_rRamAddress_2_1\ : std_logic;
signal \pEcho_rRamAddress_2_cry_0\ : std_logic;
signal \rRamAddressZ0Z_2\ : std_logic;
signal \pEcho_rRamAddress_2_2\ : std_logic;
signal \pEcho_rRamAddress_2_cry_1\ : std_logic;
signal \pEcho_rRamAddress_2_cry_2\ : std_logic;
signal \rRamAddressZ0Z_4\ : std_logic;
signal \pEcho_rRamAddress_2_4\ : std_logic;
signal \pEcho_rRamAddress_2_cry_3\ : std_logic;
signal \pEcho_rRamAddress_2_cry_4\ : std_logic;
signal \pEcho_rRamAddress_2_5\ : std_logic;
signal \pEcho_rRamAddress_2_5_cascade_\ : std_logic;
signal \rRamAddressZ0Z_5\ : std_logic;
signal \pEcho_rRamAddress_2_3\ : std_logic;
signal \rRamAddressZ0Z_3\ : std_logic;
signal \rRamReadData_0\ : std_logic;
signal \rTxByteZ0Z_4\ : std_logic;
signal \rRamReadData_1\ : std_logic;
signal \rTxByteZ0Z_5\ : std_logic;
signal \rRamReadData_2\ : std_logic;
signal \rTxByteZ0Z_6\ : std_logic;
signal \rRamReadData_3\ : std_logic;
signal \rTxByteZ0Z_7\ : std_logic;
signal \rRxReady\ : std_logic;
signal \G_11_i_a3_0_6\ : std_logic;
signal \G_11_i_a3_0_4_cascade_\ : std_logic;
signal \uartRxInst_un1_rData_0_sqmuxa_0\ : std_logic;
signal \N_5\ : std_logic;
signal \uartRxInst.un1_rCycleCounter_2_sqmuxa_0\ : std_logic;
signal \uartRxInst.rCycleCounterZ0Z_5\ : std_logic;
signal \uartRxInst.rCycleCounterZ0Z_4\ : std_logic;
signal \uartRxInst.un12_rstate_3_cascade_\ : std_logic;
signal \uartRxInst.N_83_0_i\ : std_logic;
signal \uartRxInst.N_83_0_i_cascade_\ : std_logic;
signal \uartRxInst.rState_0_sqmuxa_1_1\ : std_logic;
signal \uartRxInst.rDataCounter_0_sqmuxa\ : std_logic;
signal \uartRxInst.rCycleCounter_cry_0_THRU_CO\ : std_logic;
signal \uartRxInst.rstateZ0\ : std_logic;
signal \uartRxInst.rCycleCounter_s_2\ : std_logic;
signal \uartRxInst.un12_rstate_4\ : std_logic;
signal \uartRxInst.rCycleCounterZ0Z_1\ : std_logic;
signal \uartRxInst_rState_0\ : std_logic;
signal \uartRxInst.g0_0_5_cascade_\ : std_logic;
signal \uartRxInst.g0_0_4\ : std_logic;
signal \i_UART_RX_c\ : std_logic;
signal \uartRxInst_rState_1\ : std_logic;
signal \uartRxInst.N_83_0_i_0_cascade_\ : std_logic;
signal \uartRxInst.rCycleCounter_s_3\ : std_logic;
signal \uartRxInst.N_83_0_i_0\ : std_logic;
signal \uartRxInst.rCycleCounterZ0Z_0\ : std_logic;
signal \i_Clk_c_g\ : std_logic;
signal \uartRxInst.rCycleCountere_0_i\ : std_logic;
signal \uartRxInst.rCycleCounterZ0Z_2\ : std_logic;
signal \uartRxInst.rCycleCounterZ0Z_7\ : std_logic;
signal \uartRxInst.rCycleCounterZ0Z_3\ : std_logic;
signal \uartRxInst.rCycleCounterZ0Z_6\ : std_logic;
signal \G_11_i_a3_0_5\ : std_logic;
signal \CONSTANT_ZERO_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \i_Clk_wire\ : std_logic;
signal \o_UART_TX_wire\ : std_logic;
signal \i_UART_RX_wire\ : std_logic;
signal \ramInst.rramvalues_rramvalues_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \ramInst.rramvalues_rramvalues_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \ramInst.rramvalues_rramvalues_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \ramInst.rramvalues_rramvalues_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \ramInst.rramvalues_rramvalues_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \i_Clk_wire\ <= i_Clk;
    o_UART_TX <= \o_UART_TX_wire\;
    \i_UART_RX_wire\ <= i_UART_RX;
    \rRamReadData_3\ <= \ramInst.rramvalues_rramvalues_0_0_physical_RDATA_wire\(3);
    \rRamReadData_2\ <= \ramInst.rramvalues_rramvalues_0_0_physical_RDATA_wire\(2);
    \rRamReadData_1\ <= \ramInst.rramvalues_rramvalues_0_0_physical_RDATA_wire\(1);
    \rRamReadData_0\ <= \ramInst.rramvalues_rramvalues_0_0_physical_RDATA_wire\(0);
    \ramInst.rramvalues_rramvalues_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__2113\&\N__2134\&\N__2401\&\N__2173\&\N__2209\&\N__2236\;
    \ramInst.rramvalues_rramvalues_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__2416\&\N__2152\&\N__2386\&\N__2191\&\N__2227\&\N__2260\;
    \ramInst.rramvalues_rramvalues_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \ramInst.rramvalues_rramvalues_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';

    \ramInst.rramvalues_rramvalues_0_0_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000101100000000000011110000000000000101000000000000101000000000000000000000000000001011000000000000111100000000000000000000000000001011000000000000111100000000000001010000000000001010000000000000000000000000000010110000000000001111",
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_3 => "0000000000000000000000000000101100000000000011110000000000000101000000000000101000000000000000000000000000001011000000000000111100000000000000000000000000001011000000000000111100000000000001010000000000001010000000000000000000000000000010110000000000001111",
            INIT_2 => "0000000000000000000000000000101100000000000011110000000000000101000000000000101000000000000000000000000000001011000000000000111100000000000000000000000000001011000000000000111100000000000001010000000000001010000000000000000000000000000010110000000000001111",
            INIT_1 => "0000000000000000000000000000101100000000000011110000000000000101000000000000101000000000000000000000000000001011000000000000111100000000000000000000000000001011000000000000111100000000000001010000000000001010000000000000000000000000000010110000000000001111",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \ramInst.rramvalues_rramvalues_0_0_physical_RDATA_wire\,
            RADDR => \ramInst.rramvalues_rramvalues_0_0_physical_RADDR_wire\,
            WADDR => \ramInst.rramvalues_rramvalues_0_0_physical_WADDR_wire\,
            MASK => \ramInst.rramvalues_rramvalues_0_0_physical_MASK_wire\,
            WDATA => \ramInst.rramvalues_rramvalues_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__2789\,
            RE => \N__2009\,
            WCLKE => \N__2605\,
            WCLK => \N__2790\,
            WE => \N__2010\
        );

    \i_Clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3125\,
            GLOBALBUFFEROUTPUT => \i_Clk_c_g\
        );

    \i_Clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3127\,
            DIN => \N__3126\,
            DOUT => \N__3125\,
            PACKAGEPIN => \i_Clk_wire\
        );

    \i_Clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3127\,
            PADOUT => \N__3126\,
            PADIN => \N__3125\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_UART_TX_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3116\,
            DIN => \N__3115\,
            DOUT => \N__3114\,
            PACKAGEPIN => \o_UART_TX_wire\
        );

    \o_UART_TX_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3116\,
            PADOUT => \N__3115\,
            PADIN => \N__3114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1426\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_UART_RX_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3107\,
            DIN => \N__3106\,
            DOUT => \N__3105\,
            PACKAGEPIN => \i_UART_RX_wire\
        );

    \i_UART_RX_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3107\,
            PADOUT => \N__3106\,
            PADIN => \N__3105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \i_UART_RX_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__706\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3085\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3085\,
            I => \uartRxInst.un12_rstate_4\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__3082\,
            I => \N__3078\
        );

    \I__703\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3070\
        );

    \I__702\ : InMux
    port map (
            O => \N__3078\,
            I => \N__3070\
        );

    \I__701\ : InMux
    port map (
            O => \N__3077\,
            I => \N__3067\
        );

    \I__700\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3064\
        );

    \I__699\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3061\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3070\,
            I => \uartRxInst.rCycleCounterZ0Z_1\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3067\,
            I => \uartRxInst.rCycleCounterZ0Z_1\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3064\,
            I => \uartRxInst.rCycleCounterZ0Z_1\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3061\,
            I => \uartRxInst.rCycleCounterZ0Z_1\
        );

    \I__694\ : InMux
    port map (
            O => \N__3052\,
            I => \N__3037\
        );

    \I__693\ : InMux
    port map (
            O => \N__3051\,
            I => \N__3028\
        );

    \I__692\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3028\
        );

    \I__691\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3028\
        );

    \I__690\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3028\
        );

    \I__689\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3025\
        );

    \I__688\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3020\
        );

    \I__687\ : InMux
    port map (
            O => \N__3045\,
            I => \N__3020\
        );

    \I__686\ : InMux
    port map (
            O => \N__3044\,
            I => \N__3015\
        );

    \I__685\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3015\
        );

    \I__684\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3008\
        );

    \I__683\ : InMux
    port map (
            O => \N__3041\,
            I => \N__3008\
        );

    \I__682\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3008\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3037\,
            I => \N__3003\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3028\,
            I => \N__3003\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3025\,
            I => \uartRxInst_rState_0\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3020\,
            I => \uartRxInst_rState_0\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3015\,
            I => \uartRxInst_rState_0\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__3008\,
            I => \uartRxInst_rState_0\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__3003\,
            I => \uartRxInst_rState_0\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__2992\,
            I => \uartRxInst.g0_0_5_cascade_\
        );

    \I__673\ : InMux
    port map (
            O => \N__2989\,
            I => \N__2986\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__2986\,
            I => \uartRxInst.g0_0_4\
        );

    \I__671\ : InMux
    port map (
            O => \N__2983\,
            I => \N__2973\
        );

    \I__670\ : InMux
    port map (
            O => \N__2982\,
            I => \N__2973\
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__2981\,
            I => \N__2969\
        );

    \I__668\ : InMux
    port map (
            O => \N__2980\,
            I => \N__2964\
        );

    \I__667\ : InMux
    port map (
            O => \N__2979\,
            I => \N__2964\
        );

    \I__666\ : InMux
    port map (
            O => \N__2978\,
            I => \N__2961\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__2973\,
            I => \N__2958\
        );

    \I__664\ : InMux
    port map (
            O => \N__2972\,
            I => \N__2953\
        );

    \I__663\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2953\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__2964\,
            I => \N__2950\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__2961\,
            I => \N__2947\
        );

    \I__660\ : Span4Mux_h
    port map (
            O => \N__2958\,
            I => \N__2942\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__2953\,
            I => \N__2942\
        );

    \I__658\ : Span4Mux_v
    port map (
            O => \N__2950\,
            I => \N__2939\
        );

    \I__657\ : Span4Mux_v
    port map (
            O => \N__2947\,
            I => \N__2936\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__2942\,
            I => \N__2933\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__2939\,
            I => \i_UART_RX_c\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__2936\,
            I => \i_UART_RX_c\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__2933\,
            I => \i_UART_RX_c\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__2926\,
            I => \N__2919\
        );

    \I__651\ : InMux
    port map (
            O => \N__2925\,
            I => \N__2911\
        );

    \I__650\ : InMux
    port map (
            O => \N__2924\,
            I => \N__2911\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__2923\,
            I => \N__2905\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__2922\,
            I => \N__2902\
        );

    \I__647\ : InMux
    port map (
            O => \N__2919\,
            I => \N__2898\
        );

    \I__646\ : InMux
    port map (
            O => \N__2918\,
            I => \N__2893\
        );

    \I__645\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2893\
        );

    \I__644\ : InMux
    port map (
            O => \N__2916\,
            I => \N__2890\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__2911\,
            I => \N__2887\
        );

    \I__642\ : InMux
    port map (
            O => \N__2910\,
            I => \N__2882\
        );

    \I__641\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2882\
        );

    \I__640\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2873\
        );

    \I__639\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2873\
        );

    \I__638\ : InMux
    port map (
            O => \N__2902\,
            I => \N__2873\
        );

    \I__637\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2873\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__2898\,
            I => \uartRxInst_rState_1\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__2893\,
            I => \uartRxInst_rState_1\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__2890\,
            I => \uartRxInst_rState_1\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__2887\,
            I => \uartRxInst_rState_1\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__2882\,
            I => \uartRxInst_rState_1\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__2873\,
            I => \uartRxInst_rState_1\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__2860\,
            I => \uartRxInst.N_83_0_i_0_cascade_\
        );

    \I__629\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2854\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__2854\,
            I => \uartRxInst.rCycleCounter_s_3\
        );

    \I__627\ : InMux
    port map (
            O => \N__2851\,
            I => \N__2842\
        );

    \I__626\ : InMux
    port map (
            O => \N__2850\,
            I => \N__2835\
        );

    \I__625\ : InMux
    port map (
            O => \N__2849\,
            I => \N__2835\
        );

    \I__624\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2835\
        );

    \I__623\ : InMux
    port map (
            O => \N__2847\,
            I => \N__2828\
        );

    \I__622\ : InMux
    port map (
            O => \N__2846\,
            I => \N__2828\
        );

    \I__621\ : InMux
    port map (
            O => \N__2845\,
            I => \N__2828\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__2842\,
            I => \uartRxInst.N_83_0_i_0\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__2835\,
            I => \uartRxInst.N_83_0_i_0\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__2828\,
            I => \uartRxInst.N_83_0_i_0\
        );

    \I__617\ : InMux
    port map (
            O => \N__2821\,
            I => \N__2814\
        );

    \I__616\ : InMux
    port map (
            O => \N__2820\,
            I => \N__2811\
        );

    \I__615\ : InMux
    port map (
            O => \N__2819\,
            I => \N__2804\
        );

    \I__614\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2804\
        );

    \I__613\ : InMux
    port map (
            O => \N__2817\,
            I => \N__2804\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__2814\,
            I => \uartRxInst.rCycleCounterZ0Z_0\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__2811\,
            I => \uartRxInst.rCycleCounterZ0Z_0\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__2804\,
            I => \uartRxInst.rCycleCounterZ0Z_0\
        );

    \I__609\ : ClkMux
    port map (
            O => \N__2797\,
            I => \N__2749\
        );

    \I__608\ : ClkMux
    port map (
            O => \N__2796\,
            I => \N__2749\
        );

    \I__607\ : ClkMux
    port map (
            O => \N__2795\,
            I => \N__2749\
        );

    \I__606\ : ClkMux
    port map (
            O => \N__2794\,
            I => \N__2749\
        );

    \I__605\ : ClkMux
    port map (
            O => \N__2793\,
            I => \N__2749\
        );

    \I__604\ : ClkMux
    port map (
            O => \N__2792\,
            I => \N__2749\
        );

    \I__603\ : ClkMux
    port map (
            O => \N__2791\,
            I => \N__2749\
        );

    \I__602\ : ClkMux
    port map (
            O => \N__2790\,
            I => \N__2749\
        );

    \I__601\ : ClkMux
    port map (
            O => \N__2789\,
            I => \N__2749\
        );

    \I__600\ : ClkMux
    port map (
            O => \N__2788\,
            I => \N__2749\
        );

    \I__599\ : ClkMux
    port map (
            O => \N__2787\,
            I => \N__2749\
        );

    \I__598\ : ClkMux
    port map (
            O => \N__2786\,
            I => \N__2749\
        );

    \I__597\ : ClkMux
    port map (
            O => \N__2785\,
            I => \N__2749\
        );

    \I__596\ : ClkMux
    port map (
            O => \N__2784\,
            I => \N__2749\
        );

    \I__595\ : ClkMux
    port map (
            O => \N__2783\,
            I => \N__2749\
        );

    \I__594\ : ClkMux
    port map (
            O => \N__2782\,
            I => \N__2749\
        );

    \I__593\ : GlobalMux
    port map (
            O => \N__2749\,
            I => \N__2746\
        );

    \I__592\ : gio2CtrlBuf
    port map (
            O => \N__2746\,
            I => \i_Clk_c_g\
        );

    \I__591\ : CEMux
    port map (
            O => \N__2743\,
            I => \N__2739\
        );

    \I__590\ : CEMux
    port map (
            O => \N__2742\,
            I => \N__2736\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__2739\,
            I => \N__2732\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__2736\,
            I => \N__2729\
        );

    \I__587\ : CEMux
    port map (
            O => \N__2735\,
            I => \N__2726\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__2732\,
            I => \N__2723\
        );

    \I__585\ : Span4Mux_v
    port map (
            O => \N__2729\,
            I => \N__2720\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__2726\,
            I => \N__2717\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__2723\,
            I => \uartRxInst.rCycleCountere_0_i\
        );

    \I__582\ : Odrv4
    port map (
            O => \N__2720\,
            I => \uartRxInst.rCycleCountere_0_i\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__2717\,
            I => \uartRxInst.rCycleCountere_0_i\
        );

    \I__580\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2704\
        );

    \I__579\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2701\
        );

    \I__578\ : InMux
    port map (
            O => \N__2708\,
            I => \N__2696\
        );

    \I__577\ : InMux
    port map (
            O => \N__2707\,
            I => \N__2696\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__2704\,
            I => \uartRxInst.rCycleCounterZ0Z_2\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__2701\,
            I => \uartRxInst.rCycleCounterZ0Z_2\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__2696\,
            I => \uartRxInst.rCycleCounterZ0Z_2\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__2689\,
            I => \N__2686\
        );

    \I__572\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2680\
        );

    \I__571\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2677\
        );

    \I__570\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2674\
        );

    \I__569\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2671\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__2680\,
            I => \uartRxInst.rCycleCounterZ0Z_7\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__2677\,
            I => \uartRxInst.rCycleCounterZ0Z_7\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__2674\,
            I => \uartRxInst.rCycleCounterZ0Z_7\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__2671\,
            I => \uartRxInst.rCycleCounterZ0Z_7\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__2662\,
            I => \N__2657\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__2661\,
            I => \N__2653\
        );

    \I__562\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2650\
        );

    \I__561\ : InMux
    port map (
            O => \N__2657\,
            I => \N__2647\
        );

    \I__560\ : InMux
    port map (
            O => \N__2656\,
            I => \N__2642\
        );

    \I__559\ : InMux
    port map (
            O => \N__2653\,
            I => \N__2642\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__2650\,
            I => \uartRxInst.rCycleCounterZ0Z_3\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__2647\,
            I => \uartRxInst.rCycleCounterZ0Z_3\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__2642\,
            I => \uartRxInst.rCycleCounterZ0Z_3\
        );

    \I__555\ : InMux
    port map (
            O => \N__2635\,
            I => \N__2629\
        );

    \I__554\ : InMux
    port map (
            O => \N__2634\,
            I => \N__2626\
        );

    \I__553\ : InMux
    port map (
            O => \N__2633\,
            I => \N__2623\
        );

    \I__552\ : InMux
    port map (
            O => \N__2632\,
            I => \N__2620\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__2629\,
            I => \uartRxInst.rCycleCounterZ0Z_6\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__2626\,
            I => \uartRxInst.rCycleCounterZ0Z_6\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__2623\,
            I => \uartRxInst.rCycleCounterZ0Z_6\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2620\,
            I => \uartRxInst.rCycleCounterZ0Z_6\
        );

    \I__547\ : InMux
    port map (
            O => \N__2611\,
            I => \N__2608\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2608\,
            I => \G_11_i_a3_0_5\
        );

    \I__545\ : CEMux
    port map (
            O => \N__2605\,
            I => \N__2602\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__2602\,
            I => \N__2599\
        );

    \I__543\ : Span4Mux_v
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__2596\,
            I => \CONSTANT_ZERO_NET\
        );

    \I__541\ : InMux
    port map (
            O => \N__2593\,
            I => \N__2590\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2590\,
            I => \G_11_i_a3_0_6\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__2587\,
            I => \G_11_i_a3_0_4_cascade_\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__2584\,
            I => \N__2581\
        );

    \I__537\ : InMux
    port map (
            O => \N__2581\,
            I => \N__2577\
        );

    \I__536\ : InMux
    port map (
            O => \N__2580\,
            I => \N__2574\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__2577\,
            I => \uartRxInst_un1_rData_0_sqmuxa_0\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__2574\,
            I => \uartRxInst_un1_rData_0_sqmuxa_0\
        );

    \I__533\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2566\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__2566\,
            I => \N__2563\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__2563\,
            I => \N_5\
        );

    \I__530\ : CEMux
    port map (
            O => \N__2560\,
            I => \N__2557\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__2557\,
            I => \N__2554\
        );

    \I__528\ : Span4Mux_s3_h
    port map (
            O => \N__2554\,
            I => \N__2551\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__2551\,
            I => \uartRxInst.un1_rCycleCounter_2_sqmuxa_0\
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__2548\,
            I => \N__2541\
        );

    \I__525\ : InMux
    port map (
            O => \N__2547\,
            I => \N__2538\
        );

    \I__524\ : InMux
    port map (
            O => \N__2546\,
            I => \N__2531\
        );

    \I__523\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2531\
        );

    \I__522\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2531\
        );

    \I__521\ : InMux
    port map (
            O => \N__2541\,
            I => \N__2528\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__2538\,
            I => \uartRxInst.rCycleCounterZ0Z_5\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__2531\,
            I => \uartRxInst.rCycleCounterZ0Z_5\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__2528\,
            I => \uartRxInst.rCycleCounterZ0Z_5\
        );

    \I__517\ : InMux
    port map (
            O => \N__2521\,
            I => \N__2514\
        );

    \I__516\ : InMux
    port map (
            O => \N__2520\,
            I => \N__2509\
        );

    \I__515\ : InMux
    port map (
            O => \N__2519\,
            I => \N__2509\
        );

    \I__514\ : InMux
    port map (
            O => \N__2518\,
            I => \N__2504\
        );

    \I__513\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2504\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__2514\,
            I => \uartRxInst.rCycleCounterZ0Z_4\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__2509\,
            I => \uartRxInst.rCycleCounterZ0Z_4\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__2504\,
            I => \uartRxInst.rCycleCounterZ0Z_4\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__2497\,
            I => \uartRxInst.un12_rstate_3_cascade_\
        );

    \I__508\ : InMux
    port map (
            O => \N__2494\,
            I => \N__2488\
        );

    \I__507\ : InMux
    port map (
            O => \N__2493\,
            I => \N__2481\
        );

    \I__506\ : InMux
    port map (
            O => \N__2492\,
            I => \N__2481\
        );

    \I__505\ : InMux
    port map (
            O => \N__2491\,
            I => \N__2481\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2488\,
            I => \uartRxInst.N_83_0_i\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2481\,
            I => \uartRxInst.N_83_0_i\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__2476\,
            I => \uartRxInst.N_83_0_i_cascade_\
        );

    \I__501\ : InMux
    port map (
            O => \N__2473\,
            I => \N__2467\
        );

    \I__500\ : InMux
    port map (
            O => \N__2472\,
            I => \N__2467\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2467\,
            I => \uartRxInst.rState_0_sqmuxa_1_1\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__2464\,
            I => \N__2460\
        );

    \I__497\ : InMux
    port map (
            O => \N__2463\,
            I => \N__2452\
        );

    \I__496\ : InMux
    port map (
            O => \N__2460\,
            I => \N__2452\
        );

    \I__495\ : InMux
    port map (
            O => \N__2459\,
            I => \N__2452\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2452\,
            I => \uartRxInst.rDataCounter_0_sqmuxa\
        );

    \I__493\ : InMux
    port map (
            O => \N__2449\,
            I => \N__2446\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2446\,
            I => \uartRxInst.rCycleCounter_cry_0_THRU_CO\
        );

    \I__491\ : SRMux
    port map (
            O => \N__2443\,
            I => \N__2439\
        );

    \I__490\ : InMux
    port map (
            O => \N__2442\,
            I => \N__2436\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__2439\,
            I => \N__2433\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__2436\,
            I => \N__2430\
        );

    \I__487\ : Odrv12
    port map (
            O => \N__2433\,
            I => \uartRxInst.rstateZ0\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__2430\,
            I => \uartRxInst.rstateZ0\
        );

    \I__485\ : InMux
    port map (
            O => \N__2425\,
            I => \N__2422\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__2422\,
            I => \uartRxInst.rCycleCounter_s_2\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__2419\,
            I => \pEcho_rRamAddress_2_5_cascade_\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__2416\,
            I => \N__2413\
        );

    \I__481\ : InMux
    port map (
            O => \N__2413\,
            I => \N__2409\
        );

    \I__480\ : InMux
    port map (
            O => \N__2412\,
            I => \N__2406\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2409\,
            I => \rRamAddressZ0Z_5\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__2406\,
            I => \rRamAddressZ0Z_5\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__2401\,
            I => \N__2398\
        );

    \I__476\ : InMux
    port map (
            O => \N__2398\,
            I => \N__2394\
        );

    \I__475\ : InMux
    port map (
            O => \N__2397\,
            I => \N__2391\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2394\,
            I => \pEcho_rRamAddress_2_3\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__2391\,
            I => \pEcho_rRamAddress_2_3\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__2386\,
            I => \N__2383\
        );

    \I__471\ : InMux
    port map (
            O => \N__2383\,
            I => \N__2379\
        );

    \I__470\ : InMux
    port map (
            O => \N__2382\,
            I => \N__2376\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2379\,
            I => \rRamAddressZ0Z_3\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2376\,
            I => \rRamAddressZ0Z_3\
        );

    \I__467\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2368\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__2368\,
            I => \rRamReadData_0\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__2365\,
            I => \N__2362\
        );

    \I__464\ : InMux
    port map (
            O => \N__2362\,
            I => \N__2359\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2359\,
            I => \N__2356\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__2356\,
            I => \rTxByteZ0Z_4\
        );

    \I__461\ : InMux
    port map (
            O => \N__2353\,
            I => \N__2350\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__2350\,
            I => \rRamReadData_1\
        );

    \I__459\ : InMux
    port map (
            O => \N__2347\,
            I => \N__2344\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2344\,
            I => \rTxByteZ0Z_5\
        );

    \I__457\ : InMux
    port map (
            O => \N__2341\,
            I => \N__2338\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2338\,
            I => \rRamReadData_2\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__2335\,
            I => \N__2332\
        );

    \I__454\ : InMux
    port map (
            O => \N__2332\,
            I => \N__2329\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2329\,
            I => \N__2326\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__2326\,
            I => \rTxByteZ0Z_6\
        );

    \I__451\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2320\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2320\,
            I => \rRamReadData_3\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__2317\,
            I => \N__2314\
        );

    \I__448\ : InMux
    port map (
            O => \N__2314\,
            I => \N__2311\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2311\,
            I => \N__2308\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__2308\,
            I => \rTxByteZ0Z_7\
        );

    \I__445\ : CEMux
    port map (
            O => \N__2305\,
            I => \N__2301\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__2304\,
            I => \N__2294\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2301\,
            I => \N__2291\
        );

    \I__442\ : InMux
    port map (
            O => \N__2300\,
            I => \N__2288\
        );

    \I__441\ : InMux
    port map (
            O => \N__2299\,
            I => \N__2285\
        );

    \I__440\ : InMux
    port map (
            O => \N__2298\,
            I => \N__2282\
        );

    \I__439\ : InMux
    port map (
            O => \N__2297\,
            I => \N__2279\
        );

    \I__438\ : InMux
    port map (
            O => \N__2294\,
            I => \N__2276\
        );

    \I__437\ : Odrv4
    port map (
            O => \N__2291\,
            I => \rRxReady\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2288\,
            I => \rRxReady\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2285\,
            I => \rRxReady\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2282\,
            I => \rRxReady\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2279\,
            I => \rRxReady\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2276\,
            I => \rRxReady\
        );

    \I__431\ : InMux
    port map (
            O => \N__2263\,
            I => \uartRxInst.rCycleCounter_cry_6\
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__2260\,
            I => \N__2257\
        );

    \I__429\ : InMux
    port map (
            O => \N__2257\,
            I => \N__2254\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2254\,
            I => \N__2249\
        );

    \I__427\ : InMux
    port map (
            O => \N__2253\,
            I => \N__2246\
        );

    \I__426\ : InMux
    port map (
            O => \N__2252\,
            I => \N__2243\
        );

    \I__425\ : Odrv4
    port map (
            O => \N__2249\,
            I => \rRamAddressZ0Z_0\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__2246\,
            I => \rRamAddressZ0Z_0\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2243\,
            I => \rRamAddressZ0Z_0\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__2236\,
            I => \N__2233\
        );

    \I__421\ : InMux
    port map (
            O => \N__2233\,
            I => \N__2230\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__2230\,
            I => \pEcho_rRamAddress_2_0\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__2227\,
            I => \N__2224\
        );

    \I__418\ : InMux
    port map (
            O => \N__2224\,
            I => \N__2221\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2221\,
            I => \N__2217\
        );

    \I__416\ : InMux
    port map (
            O => \N__2220\,
            I => \N__2214\
        );

    \I__415\ : Odrv4
    port map (
            O => \N__2217\,
            I => \rRamAddressZ0Z_1\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2214\,
            I => \rRamAddressZ0Z_1\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__2209\,
            I => \N__2206\
        );

    \I__412\ : InMux
    port map (
            O => \N__2206\,
            I => \N__2202\
        );

    \I__411\ : InMux
    port map (
            O => \N__2205\,
            I => \N__2199\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2202\,
            I => \pEcho_rRamAddress_2_1\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2199\,
            I => \pEcho_rRamAddress_2_1\
        );

    \I__408\ : InMux
    port map (
            O => \N__2194\,
            I => \pEcho_rRamAddress_2_cry_0\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__2191\,
            I => \N__2188\
        );

    \I__406\ : InMux
    port map (
            O => \N__2188\,
            I => \N__2185\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2185\,
            I => \N__2181\
        );

    \I__404\ : InMux
    port map (
            O => \N__2184\,
            I => \N__2178\
        );

    \I__403\ : Odrv4
    port map (
            O => \N__2181\,
            I => \rRamAddressZ0Z_2\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2178\,
            I => \rRamAddressZ0Z_2\
        );

    \I__401\ : CascadeMux
    port map (
            O => \N__2173\,
            I => \N__2170\
        );

    \I__400\ : InMux
    port map (
            O => \N__2170\,
            I => \N__2166\
        );

    \I__399\ : InMux
    port map (
            O => \N__2169\,
            I => \N__2163\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2166\,
            I => \pEcho_rRamAddress_2_2\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2163\,
            I => \pEcho_rRamAddress_2_2\
        );

    \I__396\ : InMux
    port map (
            O => \N__2158\,
            I => \pEcho_rRamAddress_2_cry_1\
        );

    \I__395\ : InMux
    port map (
            O => \N__2155\,
            I => \pEcho_rRamAddress_2_cry_2\
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__2152\,
            I => \N__2149\
        );

    \I__393\ : InMux
    port map (
            O => \N__2149\,
            I => \N__2146\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2146\,
            I => \N__2142\
        );

    \I__391\ : InMux
    port map (
            O => \N__2145\,
            I => \N__2139\
        );

    \I__390\ : Odrv4
    port map (
            O => \N__2142\,
            I => \rRamAddressZ0Z_4\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2139\,
            I => \rRamAddressZ0Z_4\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__2134\,
            I => \N__2131\
        );

    \I__387\ : InMux
    port map (
            O => \N__2131\,
            I => \N__2127\
        );

    \I__386\ : InMux
    port map (
            O => \N__2130\,
            I => \N__2124\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2127\,
            I => \pEcho_rRamAddress_2_4\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2124\,
            I => \pEcho_rRamAddress_2_4\
        );

    \I__383\ : InMux
    port map (
            O => \N__2119\,
            I => \pEcho_rRamAddress_2_cry_3\
        );

    \I__382\ : InMux
    port map (
            O => \N__2116\,
            I => \pEcho_rRamAddress_2_cry_4\
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__2113\,
            I => \N__2110\
        );

    \I__380\ : InMux
    port map (
            O => \N__2110\,
            I => \N__2107\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2107\,
            I => \pEcho_rRamAddress_2_5\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__2104\,
            I => \N__2100\
        );

    \I__377\ : InMux
    port map (
            O => \N__2103\,
            I => \N__2096\
        );

    \I__376\ : InMux
    port map (
            O => \N__2100\,
            I => \N__2091\
        );

    \I__375\ : InMux
    port map (
            O => \N__2099\,
            I => \N__2091\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2096\,
            I => \uartRxInst.rDataCounterZ0Z_1\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2091\,
            I => \uartRxInst.rDataCounterZ0Z_1\
        );

    \I__372\ : InMux
    port map (
            O => \N__2086\,
            I => \N__2083\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2083\,
            I => \N__2077\
        );

    \I__370\ : InMux
    port map (
            O => \N__2082\,
            I => \N__2070\
        );

    \I__369\ : InMux
    port map (
            O => \N__2081\,
            I => \N__2070\
        );

    \I__368\ : InMux
    port map (
            O => \N__2080\,
            I => \N__2070\
        );

    \I__367\ : Odrv4
    port map (
            O => \N__2077\,
            I => \uartRxInst.rDataCounterZ0Z_0\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2070\,
            I => \uartRxInst.rDataCounterZ0Z_0\
        );

    \I__365\ : InMux
    port map (
            O => \N__2065\,
            I => \N__2062\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2062\,
            I => \uartRxInst.CO1_0\
        );

    \I__363\ : InMux
    port map (
            O => \N__2059\,
            I => \uartRxInst.rCycleCounter_cry_0\
        );

    \I__362\ : InMux
    port map (
            O => \N__2056\,
            I => \uartRxInst.rCycleCounter_cry_1\
        );

    \I__361\ : InMux
    port map (
            O => \N__2053\,
            I => \uartRxInst.rCycleCounter_cry_2\
        );

    \I__360\ : InMux
    port map (
            O => \N__2050\,
            I => \N__2047\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2047\,
            I => \uartRxInst.rCycleCounter_cry_3_THRU_CO\
        );

    \I__358\ : InMux
    port map (
            O => \N__2044\,
            I => \uartRxInst.rCycleCounter_cry_3\
        );

    \I__357\ : InMux
    port map (
            O => \N__2041\,
            I => \N__2038\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2038\,
            I => \uartRxInst.rCycleCounter_s_5\
        );

    \I__355\ : InMux
    port map (
            O => \N__2035\,
            I => \uartRxInst.rCycleCounter_cry_4\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__2032\,
            I => \N__2027\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__2031\,
            I => \N__2024\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__2030\,
            I => \N__2021\
        );

    \I__351\ : InMux
    port map (
            O => \N__2027\,
            I => \N__2011\
        );

    \I__350\ : InMux
    port map (
            O => \N__2024\,
            I => \N__2011\
        );

    \I__349\ : InMux
    port map (
            O => \N__2021\,
            I => \N__2011\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__2020\,
            I => \N__2006\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__2019\,
            I => \N__2003\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__2018\,
            I => \N__2000\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2011\,
            I => \N__1997\
        );

    \I__344\ : SRMux
    port map (
            O => \N__2010\,
            I => \N__1994\
        );

    \I__343\ : SRMux
    port map (
            O => \N__2009\,
            I => \N__1991\
        );

    \I__342\ : InMux
    port map (
            O => \N__2006\,
            I => \N__1984\
        );

    \I__341\ : InMux
    port map (
            O => \N__2003\,
            I => \N__1984\
        );

    \I__340\ : InMux
    port map (
            O => \N__2000\,
            I => \N__1984\
        );

    \I__339\ : Span4Mux_v
    port map (
            O => \N__1997\,
            I => \N__1979\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__1994\,
            I => \N__1979\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__1991\,
            I => \N__1976\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__1984\,
            I => \N__1973\
        );

    \I__335\ : Span4Mux_h
    port map (
            O => \N__1979\,
            I => \N__1970\
        );

    \I__334\ : Span4Mux_v
    port map (
            O => \N__1976\,
            I => \N__1967\
        );

    \I__333\ : Odrv12
    port map (
            O => \N__1973\,
            I => \CONSTANT_ONE_NET\
        );

    \I__332\ : Odrv4
    port map (
            O => \N__1970\,
            I => \CONSTANT_ONE_NET\
        );

    \I__331\ : Odrv4
    port map (
            O => \N__1967\,
            I => \CONSTANT_ONE_NET\
        );

    \I__330\ : InMux
    port map (
            O => \N__1960\,
            I => \N__1957\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__1957\,
            I => \uartRxInst.rCycleCounter_s_6\
        );

    \I__328\ : InMux
    port map (
            O => \N__1954\,
            I => \uartRxInst.rCycleCounter_cry_5\
        );

    \I__327\ : InMux
    port map (
            O => \N__1951\,
            I => \N__1943\
        );

    \I__326\ : InMux
    port map (
            O => \N__1950\,
            I => \N__1943\
        );

    \I__325\ : InMux
    port map (
            O => \N__1949\,
            I => \N__1940\
        );

    \I__324\ : InMux
    port map (
            O => \N__1948\,
            I => \N__1937\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__1943\,
            I => \uartTxInst.rBitIndexZ0Z_1\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__1940\,
            I => \uartTxInst.rBitIndexZ0Z_1\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__1937\,
            I => \uartTxInst.rBitIndexZ0Z_1\
        );

    \I__320\ : CascadeMux
    port map (
            O => \N__1930\,
            I => \N__1926\
        );

    \I__319\ : InMux
    port map (
            O => \N__1929\,
            I => \N__1923\
        );

    \I__318\ : InMux
    port map (
            O => \N__1926\,
            I => \N__1920\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__1923\,
            I => \uartTxInst.rTxByte_0_4\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1920\,
            I => \uartTxInst.rTxByte_0_4\
        );

    \I__315\ : InMux
    port map (
            O => \N__1915\,
            I => \N__1911\
        );

    \I__314\ : InMux
    port map (
            O => \N__1914\,
            I => \N__1908\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__1911\,
            I => \uartTxInst.rTxByte_0_6\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__1908\,
            I => \uartTxInst.rTxByte_0_6\
        );

    \I__311\ : InMux
    port map (
            O => \N__1903\,
            I => \N__1896\
        );

    \I__310\ : InMux
    port map (
            O => \N__1902\,
            I => \N__1893\
        );

    \I__309\ : InMux
    port map (
            O => \N__1901\,
            I => \N__1890\
        );

    \I__308\ : InMux
    port map (
            O => \N__1900\,
            I => \N__1885\
        );

    \I__307\ : InMux
    port map (
            O => \N__1899\,
            I => \N__1885\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1896\,
            I => \N__1882\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__1893\,
            I => \uartTxInst.rBitIndexZ1Z_0\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1890\,
            I => \uartTxInst.rBitIndexZ1Z_0\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__1885\,
            I => \uartTxInst.rBitIndexZ1Z_0\
        );

    \I__302\ : Odrv4
    port map (
            O => \N__1882\,
            I => \uartTxInst.rBitIndexZ1Z_0\
        );

    \I__301\ : InMux
    port map (
            O => \N__1873\,
            I => \N__1869\
        );

    \I__300\ : InMux
    port map (
            O => \N__1872\,
            I => \N__1866\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__1869\,
            I => \uartTxInst.rTxByte_0_7\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1866\,
            I => \uartTxInst.rTxByte_0_7\
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__1861\,
            I => \uartTxInst.oSerial_3_6_i_m2_ns_1_cascade_\
        );

    \I__296\ : CascadeMux
    port map (
            O => \N__1858\,
            I => \N__1855\
        );

    \I__295\ : InMux
    port map (
            O => \N__1855\,
            I => \N__1851\
        );

    \I__294\ : InMux
    port map (
            O => \N__1854\,
            I => \N__1848\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__1851\,
            I => \uartTxInst.rTxByte_0_5\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1848\,
            I => \uartTxInst.rTxByte_0_5\
        );

    \I__291\ : InMux
    port map (
            O => \N__1843\,
            I => \N__1838\
        );

    \I__290\ : InMux
    port map (
            O => \N__1842\,
            I => \N__1835\
        );

    \I__289\ : InMux
    port map (
            O => \N__1841\,
            I => \N__1832\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__1838\,
            I => \uartTxInst.rBitIndexZ0Z_2\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__1835\,
            I => \uartTxInst.rBitIndexZ0Z_2\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1832\,
            I => \uartTxInst.rBitIndexZ0Z_2\
        );

    \I__285\ : CascadeMux
    port map (
            O => \N__1825\,
            I => \uartTxInst.N_35_cascade_\
        );

    \I__284\ : InMux
    port map (
            O => \N__1822\,
            I => \N__1812\
        );

    \I__283\ : InMux
    port map (
            O => \N__1821\,
            I => \N__1809\
        );

    \I__282\ : InMux
    port map (
            O => \N__1820\,
            I => \N__1806\
        );

    \I__281\ : InMux
    port map (
            O => \N__1819\,
            I => \N__1797\
        );

    \I__280\ : InMux
    port map (
            O => \N__1818\,
            I => \N__1797\
        );

    \I__279\ : InMux
    port map (
            O => \N__1817\,
            I => \N__1797\
        );

    \I__278\ : InMux
    port map (
            O => \N__1816\,
            I => \N__1797\
        );

    \I__277\ : InMux
    port map (
            O => \N__1815\,
            I => \N__1794\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__1812\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1809\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1806\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__1797\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1794\,
            I => \uartTxInst.rTxStateZ0Z_0\
        );

    \I__271\ : InMux
    port map (
            O => \N__1783\,
            I => \N__1780\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__1780\,
            I => \uartTxInst.N_48\
        );

    \I__269\ : CascadeMux
    port map (
            O => \N__1777\,
            I => \N__1774\
        );

    \I__268\ : InMux
    port map (
            O => \N__1774\,
            I => \N__1768\
        );

    \I__267\ : InMux
    port map (
            O => \N__1773\,
            I => \N__1768\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1768\,
            I => \uartRxInst.rDataCounterZ0Z_2\
        );

    \I__265\ : CascadeMux
    port map (
            O => \N__1765\,
            I => \uartRxInst.rstateZ0_cascade_\
        );

    \I__264\ : InMux
    port map (
            O => \N__1762\,
            I => \N__1759\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1759\,
            I => \uartTxInst.N_31\
        );

    \I__262\ : CascadeMux
    port map (
            O => \N__1756\,
            I => \N__1751\
        );

    \I__261\ : CascadeMux
    port map (
            O => \N__1755\,
            I => \N__1746\
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__1754\,
            I => \N__1743\
        );

    \I__259\ : InMux
    port map (
            O => \N__1751\,
            I => \N__1734\
        );

    \I__258\ : InMux
    port map (
            O => \N__1750\,
            I => \N__1734\
        );

    \I__257\ : InMux
    port map (
            O => \N__1749\,
            I => \N__1731\
        );

    \I__256\ : InMux
    port map (
            O => \N__1746\,
            I => \N__1722\
        );

    \I__255\ : InMux
    port map (
            O => \N__1743\,
            I => \N__1722\
        );

    \I__254\ : InMux
    port map (
            O => \N__1742\,
            I => \N__1722\
        );

    \I__253\ : InMux
    port map (
            O => \N__1741\,
            I => \N__1722\
        );

    \I__252\ : InMux
    port map (
            O => \N__1740\,
            I => \N__1717\
        );

    \I__251\ : InMux
    port map (
            O => \N__1739\,
            I => \N__1717\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1734\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1731\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1722\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1717\,
            I => \uartTxInst.rTxStateZ0Z_1\
        );

    \I__246\ : InMux
    port map (
            O => \N__1708\,
            I => \N__1705\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1705\,
            I => \uartTxInst.un2_rclkcount_4\
        );

    \I__244\ : CascadeMux
    port map (
            O => \N__1702\,
            I => \uartTxInst.N_31_cascade_\
        );

    \I__243\ : InMux
    port map (
            O => \N__1699\,
            I => \N__1696\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1696\,
            I => \uartTxInst.rTxState_10_0_x2_0_o2_1_1_1\
        );

    \I__241\ : CascadeMux
    port map (
            O => \N__1693\,
            I => \uartTxInst.rTxState_10_0_x2_0_o2_1_1_1_cascade_\
        );

    \I__240\ : InMux
    port map (
            O => \N__1690\,
            I => \N__1686\
        );

    \I__239\ : InMux
    port map (
            O => \N__1689\,
            I => \N__1683\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1686\,
            I => \uartTxInst.rTxState_10_0_x2_0_o2_d_0_1\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1683\,
            I => \uartTxInst.rTxState_10_0_x2_0_o2_d_0_1\
        );

    \I__236\ : SRMux
    port map (
            O => \N__1678\,
            I => \N__1673\
        );

    \I__235\ : CascadeMux
    port map (
            O => \N__1677\,
            I => \N__1662\
        );

    \I__234\ : CascadeMux
    port map (
            O => \N__1676\,
            I => \N__1657\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1673\,
            I => \N__1653\
        );

    \I__232\ : InMux
    port map (
            O => \N__1672\,
            I => \N__1650\
        );

    \I__231\ : InMux
    port map (
            O => \N__1671\,
            I => \N__1639\
        );

    \I__230\ : InMux
    port map (
            O => \N__1670\,
            I => \N__1639\
        );

    \I__229\ : InMux
    port map (
            O => \N__1669\,
            I => \N__1639\
        );

    \I__228\ : InMux
    port map (
            O => \N__1668\,
            I => \N__1639\
        );

    \I__227\ : InMux
    port map (
            O => \N__1667\,
            I => \N__1639\
        );

    \I__226\ : InMux
    port map (
            O => \N__1666\,
            I => \N__1632\
        );

    \I__225\ : InMux
    port map (
            O => \N__1665\,
            I => \N__1632\
        );

    \I__224\ : InMux
    port map (
            O => \N__1662\,
            I => \N__1632\
        );

    \I__223\ : InMux
    port map (
            O => \N__1661\,
            I => \N__1627\
        );

    \I__222\ : InMux
    port map (
            O => \N__1660\,
            I => \N__1627\
        );

    \I__221\ : InMux
    port map (
            O => \N__1657\,
            I => \N__1622\
        );

    \I__220\ : InMux
    port map (
            O => \N__1656\,
            I => \N__1622\
        );

    \I__219\ : Odrv12
    port map (
            O => \N__1653\,
            I => \uartTxInst.rbitindex15\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1650\,
            I => \uartTxInst.rbitindex15\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1639\,
            I => \uartTxInst.rbitindex15\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__1632\,
            I => \uartTxInst.rbitindex15\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1627\,
            I => \uartTxInst.rbitindex15\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1622\,
            I => \uartTxInst.rbitindex15\
        );

    \I__213\ : InMux
    port map (
            O => \N__1609\,
            I => \N__1602\
        );

    \I__212\ : InMux
    port map (
            O => \N__1608\,
            I => \N__1593\
        );

    \I__211\ : InMux
    port map (
            O => \N__1607\,
            I => \N__1593\
        );

    \I__210\ : InMux
    port map (
            O => \N__1606\,
            I => \N__1593\
        );

    \I__209\ : InMux
    port map (
            O => \N__1605\,
            I => \N__1593\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1602\,
            I => \N__1590\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1593\,
            I => \rTxDVZ0\
        );

    \I__206\ : Odrv4
    port map (
            O => \N__1590\,
            I => \rTxDVZ0\
        );

    \I__205\ : CascadeMux
    port map (
            O => \N__1585\,
            I => \uartRxInst.rDataCounter_RNO_0Z0Z_1_cascade_\
        );

    \I__204\ : CascadeMux
    port map (
            O => \N__1582\,
            I => \uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_\
        );

    \I__203\ : InMux
    port map (
            O => \N__1579\,
            I => \N__1574\
        );

    \I__202\ : InMux
    port map (
            O => \N__1578\,
            I => \N__1571\
        );

    \I__201\ : InMux
    port map (
            O => \N__1577\,
            I => \N__1568\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1574\,
            I => \uartTxInst.rClkCountZ0Z_6\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1571\,
            I => \uartTxInst.rClkCountZ0Z_6\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1568\,
            I => \uartTxInst.rClkCountZ0Z_6\
        );

    \I__197\ : CascadeMux
    port map (
            O => \N__1561\,
            I => \N__1557\
        );

    \I__196\ : InMux
    port map (
            O => \N__1560\,
            I => \N__1552\
        );

    \I__195\ : InMux
    port map (
            O => \N__1557\,
            I => \N__1547\
        );

    \I__194\ : InMux
    port map (
            O => \N__1556\,
            I => \N__1547\
        );

    \I__193\ : InMux
    port map (
            O => \N__1555\,
            I => \N__1544\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__1552\,
            I => \uartTxInst.rClkCountZ0Z_5\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1547\,
            I => \uartTxInst.rClkCountZ0Z_5\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1544\,
            I => \uartTxInst.rClkCountZ0Z_5\
        );

    \I__189\ : CascadeMux
    port map (
            O => \N__1537\,
            I => \N__1532\
        );

    \I__188\ : InMux
    port map (
            O => \N__1536\,
            I => \N__1525\
        );

    \I__187\ : InMux
    port map (
            O => \N__1535\,
            I => \N__1525\
        );

    \I__186\ : InMux
    port map (
            O => \N__1532\,
            I => \N__1525\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__1525\,
            I => \uartTxInst.un5_rclkcount_c4\
        );

    \I__184\ : InMux
    port map (
            O => \N__1522\,
            I => \N__1508\
        );

    \I__183\ : InMux
    port map (
            O => \N__1521\,
            I => \N__1508\
        );

    \I__182\ : InMux
    port map (
            O => \N__1520\,
            I => \N__1505\
        );

    \I__181\ : InMux
    port map (
            O => \N__1519\,
            I => \N__1500\
        );

    \I__180\ : InMux
    port map (
            O => \N__1518\,
            I => \N__1500\
        );

    \I__179\ : InMux
    port map (
            O => \N__1517\,
            I => \N__1497\
        );

    \I__178\ : InMux
    port map (
            O => \N__1516\,
            I => \N__1494\
        );

    \I__177\ : InMux
    port map (
            O => \N__1515\,
            I => \N__1487\
        );

    \I__176\ : InMux
    port map (
            O => \N__1514\,
            I => \N__1487\
        );

    \I__175\ : InMux
    port map (
            O => \N__1513\,
            I => \N__1487\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1508\,
            I => \N__1484\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1505\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1500\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__171\ : LocalMux
    port map (
            O => \N__1497\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1494\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__169\ : LocalMux
    port map (
            O => \N__1487\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__168\ : Odrv4
    port map (
            O => \N__1484\,
            I => \uartTxInst.SUM_N_3_mux\
        );

    \I__167\ : CascadeMux
    port map (
            O => \N__1471\,
            I => \N__1468\
        );

    \I__166\ : InMux
    port map (
            O => \N__1468\,
            I => \N__1461\
        );

    \I__165\ : InMux
    port map (
            O => \N__1467\,
            I => \N__1458\
        );

    \I__164\ : InMux
    port map (
            O => \N__1466\,
            I => \N__1451\
        );

    \I__163\ : InMux
    port map (
            O => \N__1465\,
            I => \N__1451\
        );

    \I__162\ : InMux
    port map (
            O => \N__1464\,
            I => \N__1451\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1461\,
            I => \N__1448\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1458\,
            I => \uartTxInst.rClkCountZ0Z_4\
        );

    \I__159\ : LocalMux
    port map (
            O => \N__1451\,
            I => \uartTxInst.rClkCountZ0Z_4\
        );

    \I__158\ : Odrv4
    port map (
            O => \N__1448\,
            I => \uartTxInst.rClkCountZ0Z_4\
        );

    \I__157\ : CascadeMux
    port map (
            O => \N__1441\,
            I => \uartTxInst.g2_0_cascade_\
        );

    \I__156\ : CascadeMux
    port map (
            O => \N__1438\,
            I => \uartTxInst.rBitIndex_RNO_0Z0Z_1_cascade_\
        );

    \I__155\ : InMux
    port map (
            O => \N__1435\,
            I => \N__1432\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1432\,
            I => \uartTxInst.rTxByte_0_sqmuxa\
        );

    \I__153\ : CascadeMux
    port map (
            O => \N__1429\,
            I => \uartTxInst.rTxState_10_0_i_a2_1_2_0_cascade_\
        );

    \I__152\ : IoInMux
    port map (
            O => \N__1426\,
            I => \N__1423\
        );

    \I__151\ : LocalMux
    port map (
            O => \N__1423\,
            I => \N__1420\
        );

    \I__150\ : IoSpan4Mux
    port map (
            O => \N__1420\,
            I => \N__1416\
        );

    \I__149\ : CascadeMux
    port map (
            O => \N__1419\,
            I => \N__1413\
        );

    \I__148\ : Span4Mux_s2_h
    port map (
            O => \N__1416\,
            I => \N__1410\
        );

    \I__147\ : InMux
    port map (
            O => \N__1413\,
            I => \N__1407\
        );

    \I__146\ : Odrv4
    port map (
            O => \N__1410\,
            I => \o_UART_TX_c\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__1407\,
            I => \o_UART_TX_c\
        );

    \I__144\ : CascadeMux
    port map (
            O => \N__1402\,
            I => \uartTxInst.rbitindex15_cascade_\
        );

    \I__143\ : InMux
    port map (
            O => \N__1399\,
            I => \N__1388\
        );

    \I__142\ : InMux
    port map (
            O => \N__1398\,
            I => \N__1388\
        );

    \I__141\ : InMux
    port map (
            O => \N__1397\,
            I => \N__1388\
        );

    \I__140\ : InMux
    port map (
            O => \N__1396\,
            I => \N__1383\
        );

    \I__139\ : InMux
    port map (
            O => \N__1395\,
            I => \N__1383\
        );

    \I__138\ : LocalMux
    port map (
            O => \N__1388\,
            I => \uartTxInst.rClkCountZ0Z_1\
        );

    \I__137\ : LocalMux
    port map (
            O => \N__1383\,
            I => \uartTxInst.rClkCountZ0Z_1\
        );

    \I__136\ : CascadeMux
    port map (
            O => \N__1378\,
            I => \uartTxInst.un2_rclkcount_5_0_cascade_\
        );

    \I__135\ : InMux
    port map (
            O => \N__1375\,
            I => \N__1371\
        );

    \I__134\ : InMux
    port map (
            O => \N__1374\,
            I => \N__1368\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__1371\,
            I => \uartTxInst.rClkCountZ0Z_7\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__1368\,
            I => \uartTxInst.rClkCountZ0Z_7\
        );

    \I__131\ : InMux
    port map (
            O => \N__1363\,
            I => \N__1356\
        );

    \I__130\ : InMux
    port map (
            O => \N__1362\,
            I => \N__1356\
        );

    \I__129\ : InMux
    port map (
            O => \N__1361\,
            I => \N__1353\
        );

    \I__128\ : LocalMux
    port map (
            O => \N__1356\,
            I => \uartTxInst.rClkCountZ0Z_3\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1353\,
            I => \uartTxInst.rClkCountZ0Z_3\
        );

    \I__126\ : CascadeMux
    port map (
            O => \N__1348\,
            I => \N__1343\
        );

    \I__125\ : CascadeMux
    port map (
            O => \N__1347\,
            I => \N__1340\
        );

    \I__124\ : InMux
    port map (
            O => \N__1346\,
            I => \N__1331\
        );

    \I__123\ : InMux
    port map (
            O => \N__1343\,
            I => \N__1331\
        );

    \I__122\ : InMux
    port map (
            O => \N__1340\,
            I => \N__1331\
        );

    \I__121\ : InMux
    port map (
            O => \N__1339\,
            I => \N__1326\
        );

    \I__120\ : InMux
    port map (
            O => \N__1338\,
            I => \N__1326\
        );

    \I__119\ : LocalMux
    port map (
            O => \N__1331\,
            I => \uartTxInst.rClkCountZ0Z_2\
        );

    \I__118\ : LocalMux
    port map (
            O => \N__1326\,
            I => \uartTxInst.rClkCountZ0Z_2\
        );

    \I__117\ : InMux
    port map (
            O => \N__1321\,
            I => \N__1306\
        );

    \I__116\ : InMux
    port map (
            O => \N__1320\,
            I => \N__1306\
        );

    \I__115\ : InMux
    port map (
            O => \N__1319\,
            I => \N__1306\
        );

    \I__114\ : InMux
    port map (
            O => \N__1318\,
            I => \N__1306\
        );

    \I__113\ : InMux
    port map (
            O => \N__1317\,
            I => \N__1299\
        );

    \I__112\ : InMux
    port map (
            O => \N__1316\,
            I => \N__1299\
        );

    \I__111\ : InMux
    port map (
            O => \N__1315\,
            I => \N__1299\
        );

    \I__110\ : LocalMux
    port map (
            O => \N__1306\,
            I => \uartTxInst.rClkCountZ0Z_0\
        );

    \I__109\ : LocalMux
    port map (
            O => \N__1299\,
            I => \uartTxInst.rClkCountZ0Z_0\
        );

    \I__108\ : CascadeMux
    port map (
            O => \N__1294\,
            I => \uartTxInst.un2_rclkcount_4_cascade_\
        );

    \I__107\ : InMux
    port map (
            O => \N__1291\,
            I => \N__1288\
        );

    \I__106\ : LocalMux
    port map (
            O => \N__1288\,
            I => \uartTxInst.un2_rclkcount_5_0\
        );

    \I__105\ : CascadeMux
    port map (
            O => \N__1285\,
            I => \uartTxInst.un5_rclkcount_c4_cascade_\
        );

    \I__104\ : CascadeMux
    port map (
            O => \N__1282\,
            I => \uartTxInst.un5_rclkcount_ac0_11_cascade_\
        );

    \I__103\ : CascadeMux
    port map (
            O => \N__1279\,
            I => \uartTxInst.un5_rclkcount_c3_cascade_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNIA4KC_3_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1318\,
            in1 => \N__1397\,
            in2 => \N__1347\,
            in3 => \N__1362\,
            lcout => \uartTxInst.un5_rclkcount_c4\,
            ltout => \uartTxInst.un5_rclkcount_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNO_0_7_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1579\,
            in1 => \N__1560\,
            in2 => \N__1285\,
            in3 => \N__1467\,
            lcout => OPEN,
            ltout => \uartTxInst.un5_rclkcount_ac0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_7_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__1661\,
            in1 => \N__1375\,
            in2 => \N__1282\,
            in3 => \N__1519\,
            lcout => \uartTxInst.rClkCountZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__1399\,
            in1 => \N__1346\,
            in2 => \N__1676\,
            in3 => \N__1320\,
            lcout => \uartTxInst.rClkCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNO_0_3_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__1319\,
            in1 => \N__1398\,
            in2 => \N__1348\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \uartTxInst.un5_rclkcount_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_3_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__1363\,
            in1 => \N__1660\,
            in2 => \N__1279\,
            in3 => \N__1516\,
            lcout => \uartTxInst.rClkCountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_0_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__1321\,
            in1 => \N__1656\,
            in2 => \_gnd_net_\,
            in3 => \N__1518\,
            lcout => \uartTxInst.rClkCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxState_RNINSDP_0_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__1820\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1739\,
            lcout => \uartTxInst.rbitindex15\,
            ltout => \uartTxInst.rbitindex15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1317\,
            in2 => \N__1402\,
            in3 => \N__1396\,
            lcout => \uartTxInst.rClkCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNI85A6_5_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1395\,
            in2 => \_gnd_net_\,
            in3 => \N__1555\,
            lcout => \uartTxInst.un2_rclkcount_5_0\,
            ltout => \uartTxInst.un2_rclkcount_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNI85BP_2_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__1316\,
            in1 => \N__1740\,
            in2 => \N__1378\,
            in3 => \N__1339\,
            lcout => \uartTxInst.rTxState_10_0_x2_0_o2_d_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxDV_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2300\,
            lcout => \rTxDVZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNIOIKC_7_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1374\,
            in1 => \N__1577\,
            in2 => \N__1471\,
            in3 => \N__1361\,
            lcout => \uartTxInst.un2_rclkcount_4\,
            ltout => \uartTxInst.un2_rclkcount_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNI4P8P_2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__1338\,
            in1 => \N__1315\,
            in2 => \N__1294\,
            in3 => \N__1291\,
            lcout => \uartTxInst.SUM_N_3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxState_1_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__1818\,
            in1 => \_gnd_net_\,
            in2 => \N__1755\,
            in3 => \N__1515\,
            lcout => \uartTxInst.rTxStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNO_1_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1816\,
            in2 => \_gnd_net_\,
            in3 => \N__1901\,
            lcout => OPEN,
            ltout => \uartTxInst.g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNO_0_1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110010"
        )
    port map (
            in0 => \N__1742\,
            in1 => \N__1513\,
            in2 => \N__1441\,
            in3 => \N__1950\,
            lcout => OPEN,
            ltout => \uartTxInst.rBitIndex_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__1690\,
            in1 => \N__1672\,
            in2 => \N__1438\,
            in3 => \N__1699\,
            lcout => \uartTxInst.rBitIndexZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxState_RNO_1_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__1609\,
            in1 => \N__1741\,
            in2 => \_gnd_net_\,
            in3 => \N__1817\,
            lcout => \uartTxInst.rTxByte_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxState_RNO_0_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__1762\,
            in1 => \N__1842\,
            in2 => \N__1754\,
            in3 => \N__1951\,
            lcout => OPEN,
            ltout => \uartTxInst.rTxState_10_0_i_a2_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxState_0_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111101100"
        )
    port map (
            in0 => \N__1514\,
            in1 => \N__1435\,
            in2 => \N__1429\,
            in3 => \N__1819\,
            lcout => \uartTxInst.rTxStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.oSerial_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__1521\,
            in1 => \N__1750\,
            in2 => \N__1419\,
            in3 => \N__1783\,
            lcout => \o_UART_TX_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => 'H',
            sr => \N__1678\
        );

    \uartTxInst.rBitIndex_0_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101001000101"
        )
    port map (
            in0 => \N__1822\,
            in1 => \N__1522\,
            in2 => \N__1756\,
            in3 => \N__1902\,
            lcout => \uartTxInst.rBitIndexZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => 'H',
            sr => \N__1678\
        );

    \CONSTANT_ONE_LUT4_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_RNO_0_6_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__1578\,
            in1 => \N__1556\,
            in2 => \N__1537\,
            in3 => \N__1464\,
            lcout => OPEN,
            ltout => \uartTxInst.rClkCount_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_6_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1517\,
            in2 => \N__1582\,
            in3 => \N__1666\,
            lcout => \uartTxInst.rClkCountZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRamAddress_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__2299\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2253\,
            lcout => \rRamAddressZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_5_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__1465\,
            in1 => \N__1665\,
            in2 => \N__1561\,
            in3 => \N__1536\,
            lcout => \uartTxInst.rClkCountZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRamAddress_2_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2169\,
            lcout => \rRamAddressZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRamAddress_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2205\,
            lcout => \rRamAddressZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rClkCount_4_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__1535\,
            in1 => \N__1466\,
            in2 => \N__1677\,
            in3 => \N__1520\,
            lcout => \uartTxInst.rClkCountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2785\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxByte_7_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__1671\,
            in1 => \N__1608\,
            in2 => \N__2317\,
            in3 => \N__1873\,
            lcout => \uartTxInst.rTxByte_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxByte_4_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__1605\,
            in1 => \N__1668\,
            in2 => \N__2365\,
            in3 => \N__1929\,
            lcout => \uartTxInst.rTxByte_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxByte_6_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__1670\,
            in1 => \N__1607\,
            in2 => \N__2335\,
            in3 => \N__1915\,
            lcout => \uartTxInst.rTxByte_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNI0NON_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1815\,
            in2 => \_gnd_net_\,
            in3 => \N__1903\,
            lcout => \uartTxInst.N_31\,
            ltout => \uartTxInst.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_RNIQ26S1_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111111"
        )
    port map (
            in0 => \N__1749\,
            in1 => \N__1708\,
            in2 => \N__1702\,
            in3 => \N__1949\,
            lcout => \uartTxInst.rTxState_10_0_x2_0_o2_1_1_1\,
            ltout => \uartTxInst.rTxState_10_0_x2_0_o2_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rBitIndex_2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100001"
        )
    port map (
            in0 => \N__1843\,
            in1 => \N__1667\,
            in2 => \N__1693\,
            in3 => \N__1689\,
            lcout => \uartTxInst.rBitIndexZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.rTxByte_5_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__1669\,
            in1 => \N__1606\,
            in2 => \N__1858\,
            in3 => \N__2347\,
            lcout => \uartTxInst.rTxByte_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rDataReady_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__2916\,
            in1 => \N__3047\,
            in2 => \_gnd_net_\,
            in3 => \N__2298\,
            lcout => \rRxReady\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rDataCounter_RNO_0_1_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001011110000"
        )
    port map (
            in0 => \N__2081\,
            in1 => \N__3043\,
            in2 => \N__2104\,
            in3 => \N__2491\,
            lcout => OPEN,
            ltout => \uartRxInst.rDataCounter_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rDataCounter_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1585\,
            in3 => \N__2459\,
            lcout => \uartRxInst.rDataCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2792\,
            ce => 'H',
            sr => \N__2443\
        );

    \uartRxInst.rDataCounter_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100111111010"
        )
    port map (
            in0 => \N__2082\,
            in1 => \N__3044\,
            in2 => \N__2464\,
            in3 => \N__2492\,
            lcout => \uartRxInst.rDataCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2792\,
            ce => 'H',
            sr => \N__2443\
        );

    \uartRxInst.rDataCounter_RNILM1D1_2_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__1773\,
            in1 => \N__2099\,
            in2 => \_gnd_net_\,
            in3 => \N__2080\,
            lcout => \uartRxInst.rState_0_sqmuxa_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.oSerial_RNO_2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__1948\,
            in1 => \N__1899\,
            in2 => \N__1930\,
            in3 => \N__1914\,
            lcout => OPEN,
            ltout => \uartTxInst.oSerial_3_6_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.oSerial_RNO_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__1900\,
            in1 => \N__1872\,
            in2 => \N__1861\,
            in3 => \N__1854\,
            lcout => OPEN,
            ltout => \uartTxInst.N_35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartTxInst.oSerial_RNO_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1841\,
            in2 => \N__1825\,
            in3 => \N__1821\,
            lcout => \uartTxInst.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rDataCounter_2_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101111000"
        )
    port map (
            in0 => \N__2493\,
            in1 => \N__2065\,
            in2 => \N__1777\,
            in3 => \N__2463\,
            lcout => \uartRxInst.rDataCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2792\,
            ce => 'H',
            sr => \N__2443\
        );

    \uartRxInst.rCycleCounter_RNI66KJ1_7_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2517\,
            in1 => \N__2684\,
            in2 => \N__2548\,
            in3 => \N__2633\,
            lcout => \uartRxInst.g0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rState_RNIRJB_0_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__3041\,
            in1 => \N__2910\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uartRxInst.rstateZ0\,
            ltout => \uartRxInst.rstateZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_5_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__2979\,
            in1 => \N__2848\,
            in2 => \N__1765\,
            in3 => \N__2041\,
            lcout => \uartRxInst.rCycleCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2794\,
            ce => \N__2735\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_6_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__2849\,
            in1 => \N__2980\,
            in2 => \N__2926\,
            in3 => \N__1960\,
            lcout => \uartRxInst.rCycleCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2794\,
            ce => \N__2735\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rState_RNIRJB_1_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__3042\,
            in1 => \N__2909\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uartRxInst.rCycleCountere_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_4_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000011101"
        )
    port map (
            in0 => \N__2518\,
            in1 => \N__2850\,
            in2 => \N__2584\,
            in3 => \N__2050\,
            lcout => \uartRxInst.rCycleCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2794\,
            ce => \N__2735\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rDataCounter_RNO_0_2_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__3040\,
            in1 => \N__2103\,
            in2 => \_gnd_net_\,
            in3 => \N__2086\,
            lcout => \uartRxInst.CO1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_cry_c_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2820\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \uartRxInst.rCycleCounter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_cry_0_THRU_LUT4_0_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3077\,
            in2 => \N__2020\,
            in3 => \N__2059\,
            lcout => \uartRxInst.rCycleCounter_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \uartRxInst.rCycleCounter_cry_0\,
            carryout => \uartRxInst.rCycleCounter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNO_0_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2709\,
            in2 => \N__2030\,
            in3 => \N__2056\,
            lcout => \uartRxInst.rCycleCounter_s_2\,
            ltout => OPEN,
            carryin => \uartRxInst.rCycleCounter_cry_1\,
            carryout => \uartRxInst.rCycleCounter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNO_0_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2660\,
            in2 => \N__2018\,
            in3 => \N__2053\,
            lcout => \uartRxInst.rCycleCounter_s_3\,
            ltout => OPEN,
            carryin => \uartRxInst.rCycleCounter_cry_2\,
            carryout => \uartRxInst.rCycleCounter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_cry_3_THRU_LUT4_0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2521\,
            in2 => \N__2032\,
            in3 => \N__2044\,
            lcout => \uartRxInst.rCycleCounter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \uartRxInst.rCycleCounter_cry_3\,
            carryout => \uartRxInst.rCycleCounter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNO_0_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2547\,
            in2 => \N__2019\,
            in3 => \N__2035\,
            lcout => \uartRxInst.rCycleCounter_s_5\,
            ltout => OPEN,
            carryin => \uartRxInst.rCycleCounter_cry_4\,
            carryout => \uartRxInst.rCycleCounter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNO_0_6_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2635\,
            in2 => \N__2031\,
            in3 => \N__1954\,
            lcout => \uartRxInst.rCycleCounter_s_6\,
            ltout => OPEN,
            carryin => \uartRxInst.rCycleCounter_cry_5\,
            carryout => \uartRxInst.rCycleCounter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_7_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010001000111"
        )
    port map (
            in0 => \N__2580\,
            in1 => \N__2851\,
            in2 => \N__2689\,
            in3 => \N__2263\,
            lcout => \uartRxInst.rCycleCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2796\,
            ce => \N__2742\,
            sr => \_gnd_net_\
        );

    \rRamAddress_4_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2130\,
            lcout => \rRamAddressZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRamAddress_RNIJ99L_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2252\,
            in2 => \N__2304\,
            in3 => \N__2297\,
            lcout => \pEcho_rRamAddress_2_0\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \pEcho_rRamAddress_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pEcho_rRamAddress_2_cry_0_c_RNI5QRQ_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2220\,
            in2 => \_gnd_net_\,
            in3 => \N__2194\,
            lcout => \pEcho_rRamAddress_2_1\,
            ltout => OPEN,
            carryin => \pEcho_rRamAddress_2_cry_0\,
            carryout => \pEcho_rRamAddress_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pEcho_rRamAddress_2_cry_1_c_RNI7TSQ_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2184\,
            in2 => \_gnd_net_\,
            in3 => \N__2158\,
            lcout => \pEcho_rRamAddress_2_2\,
            ltout => OPEN,
            carryin => \pEcho_rRamAddress_2_cry_1\,
            carryout => \pEcho_rRamAddress_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pEcho_rRamAddress_2_cry_2_c_RNI90UQ_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2382\,
            in2 => \_gnd_net_\,
            in3 => \N__2155\,
            lcout => \pEcho_rRamAddress_2_3\,
            ltout => OPEN,
            carryin => \pEcho_rRamAddress_2_cry_2\,
            carryout => \pEcho_rRamAddress_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pEcho_rRamAddress_2_cry_3_c_RNIB3VQ_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2145\,
            in2 => \_gnd_net_\,
            in3 => \N__2119\,
            lcout => \pEcho_rRamAddress_2_4\,
            ltout => OPEN,
            carryin => \pEcho_rRamAddress_2_cry_3\,
            carryout => \pEcho_rRamAddress_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pEcho_rRamAddress_2_cry_4_c_RNID60R_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2412\,
            in2 => \_gnd_net_\,
            in3 => \N__2116\,
            lcout => \pEcho_rRamAddress_2_5\,
            ltout => \pEcho_rRamAddress_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRamAddress_5_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2419\,
            in3 => \_gnd_net_\,
            lcout => \rRamAddressZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRamAddress_3_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2397\,
            lcout => \rRamAddressZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_e_0_4_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2371\,
            lcout => \rTxByteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2305\,
            sr => \_gnd_net_\
        );

    \rTxByte_e_0_5_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2353\,
            lcout => \rTxByteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2305\,
            sr => \_gnd_net_\
        );

    \rTxByte_e_0_6_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2341\,
            lcout => \rTxByteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2305\,
            sr => \_gnd_net_\
        );

    \rTxByte_e_0_7_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2323\,
            lcout => \rTxByteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2305\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rState_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111001100"
        )
    port map (
            in0 => \N__2983\,
            in1 => \N__2918\,
            in2 => \_gnd_net_\,
            in3 => \N__3046\,
            lcout => \uartRxInst_rState_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2795\,
            ce => \N__2560\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rState_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__2982\,
            in1 => \N__2917\,
            in2 => \_gnd_net_\,
            in3 => \N__3045\,
            lcout => \uartRxInst_rState_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2795\,
            ce => \N__2560\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNICOS61_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__2545\,
            in1 => \N__2520\,
            in2 => \N__2922\,
            in3 => \N__3076\,
            lcout => \G_11_i_a3_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNIAMVP_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3048\,
            in1 => \N__2544\,
            in2 => \_gnd_net_\,
            in3 => \N__2821\,
            lcout => OPEN,
            ltout => \G_11_i_a3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i_UART_RX_ibuf_RNI5MUN3_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__2569\,
            in1 => \N__2593\,
            in2 => \N__2587\,
            in3 => \N__2611\,
            lcout => \uartRxInst_un1_rData_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i_UART_RX_ibuf_RNID5E3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3049\,
            in1 => \N__2901\,
            in2 => \_gnd_net_\,
            in3 => \N__2978\,
            lcout => \N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rState_RNIC6LK4_1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111000011"
        )
    port map (
            in0 => \N__2473\,
            in1 => \N__3051\,
            in2 => \N__2923\,
            in3 => \N__2494\,
            lcout => \uartRxInst.un1_rCycleCounter_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNI55QP_7_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__2683\,
            in1 => \N__2632\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \uartRxInst.un12_rstate_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNISR773_4_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2546\,
            in1 => \N__2519\,
            in2 => \N__2497\,
            in3 => \N__3088\,
            lcout => \uartRxInst.N_83_0_i\,
            ltout => \uartRxInst.N_83_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rState_RNIC6LK4_0_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3050\,
            in1 => \N__2908\,
            in2 => \N__2476\,
            in3 => \N__2472\,
            lcout => \uartRxInst.rDataCounter_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2847\,
            in1 => \N__2449\,
            in2 => \_gnd_net_\,
            in3 => \N__3081\,
            lcout => \uartRxInst.rCycleCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2797\,
            ce => \N__2743\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_2_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__2442\,
            in1 => \N__2425\,
            in2 => \N__2981\,
            in3 => \N__2845\,
            lcout => \uartRxInst.rCycleCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2797\,
            ce => \N__2743\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNIMLJJ1_0_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3075\,
            in1 => \N__2817\,
            in2 => \N__2661\,
            in3 => \N__2707\,
            lcout => \uartRxInst.un12_rstate_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNIMLJJ1_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2818\,
            in1 => \N__2656\,
            in2 => \N__3082\,
            in3 => \N__2710\,
            lcout => OPEN,
            ltout => \uartRxInst.g0_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rState_RNINFJ73_1_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100010001"
        )
    port map (
            in0 => \N__2924\,
            in1 => \N__3052\,
            in2 => \N__2992\,
            in3 => \N__2989\,
            lcout => \uartRxInst.N_83_0_i_0\,
            ltout => \uartRxInst.N_83_0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111111010000"
        )
    port map (
            in0 => \N__2972\,
            in1 => \N__2925\,
            in2 => \N__2860\,
            in3 => \N__2857\,
            lcout => \uartRxInst.rCycleCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2797\,
            ce => \N__2743\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_0_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2846\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2819\,
            lcout => \uartRxInst.rCycleCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2797\,
            ce => \N__2743\,
            sr => \_gnd_net_\
        );

    \uartRxInst.rCycleCounter_RNI22KJ1_7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2708\,
            in1 => \N__2685\,
            in2 => \N__2662\,
            in3 => \N__2634\,
            lcout => \G_11_i_a3_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ZERO_LUT4_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ZERO_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
