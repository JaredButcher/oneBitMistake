-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 28 2019 23:31:20

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "uartRx" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of uartRx
entity uartRx is
port (
    oData : out std_logic_vector(7 downto 0);
    iClk : in std_logic;
    oDataReady : out std_logic;
    iSerial : in std_logic);
end uartRx;

-- Architecture of uartRx
-- View name is \INTERFACE\
architecture \INTERFACE\ of uartRx is

signal \N__2412\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2182\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2078\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2068\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2066\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2061\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2053\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2005\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1987\ : std_logic;
signal \N__1986\ : std_logic;
signal \N__1983\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1978\ : std_logic;
signal \N__1975\ : std_logic;
signal \N__1974\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1969\ : std_logic;
signal \N__1968\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1944\ : std_logic;
signal \N__1941\ : std_logic;
signal \N__1938\ : std_logic;
signal \N__1935\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1929\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1912\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1902\ : std_logic;
signal \N__1899\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1889\ : std_logic;
signal \N__1886\ : std_logic;
signal \N__1881\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1853\ : std_logic;
signal \N__1850\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1839\ : std_logic;
signal \N__1836\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1830\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1827\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1824\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1821\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1818\ : std_logic;
signal \N__1785\ : std_logic;
signal \N__1782\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1776\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1767\ : std_logic;
signal \N__1766\ : std_logic;
signal \N__1761\ : std_logic;
signal \N__1760\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1758\ : std_logic;
signal \N__1757\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1753\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1741\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1728\ : std_logic;
signal \N__1725\ : std_logic;
signal \N__1722\ : std_logic;
signal \N__1719\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1716\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1700\ : std_logic;
signal \N__1695\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1691\ : std_logic;
signal \N__1690\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1679\ : std_logic;
signal \N__1676\ : std_logic;
signal \N__1673\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1652\ : std_logic;
signal \N__1649\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1640\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1631\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1614\ : std_logic;
signal \N__1613\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1611\ : std_logic;
signal \N__1608\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1595\ : std_logic;
signal \N__1594\ : std_logic;
signal \N__1591\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1577\ : std_logic;
signal \N__1572\ : std_logic;
signal \N__1563\ : std_logic;
signal \N__1562\ : std_logic;
signal \N__1559\ : std_logic;
signal \N__1558\ : std_logic;
signal \N__1557\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1542\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1539\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1521\ : std_logic;
signal \N__1512\ : std_logic;
signal \N__1509\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1504\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1501\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1498\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1482\ : std_logic;
signal \N__1473\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1462\ : std_logic;
signal \N__1459\ : std_logic;
signal \N__1456\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1450\ : std_logic;
signal \N__1449\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1447\ : std_logic;
signal \N__1446\ : std_logic;
signal \N__1445\ : std_logic;
signal \N__1444\ : std_logic;
signal \N__1443\ : std_logic;
signal \N__1440\ : std_logic;
signal \N__1437\ : std_logic;
signal \N__1434\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1402\ : std_logic;
signal \N__1399\ : std_logic;
signal \N__1398\ : std_logic;
signal \N__1397\ : std_logic;
signal \N__1394\ : std_logic;
signal \N__1391\ : std_logic;
signal \N__1390\ : std_logic;
signal \N__1389\ : std_logic;
signal \N__1386\ : std_logic;
signal \N__1383\ : std_logic;
signal \N__1382\ : std_logic;
signal \N__1379\ : std_logic;
signal \N__1374\ : std_logic;
signal \N__1369\ : std_logic;
signal \N__1368\ : std_logic;
signal \N__1363\ : std_logic;
signal \N__1360\ : std_logic;
signal \N__1357\ : std_logic;
signal \N__1352\ : std_logic;
signal \N__1349\ : std_logic;
signal \N__1346\ : std_logic;
signal \N__1335\ : std_logic;
signal \N__1332\ : std_logic;
signal \N__1329\ : std_logic;
signal \N__1326\ : std_logic;
signal \N__1323\ : std_logic;
signal \N__1320\ : std_logic;
signal \N__1317\ : std_logic;
signal \N__1314\ : std_logic;
signal \N__1311\ : std_logic;
signal \N__1308\ : std_logic;
signal \N__1307\ : std_logic;
signal \N__1306\ : std_logic;
signal \N__1305\ : std_logic;
signal \N__1304\ : std_logic;
signal \N__1301\ : std_logic;
signal \N__1298\ : std_logic;
signal \N__1295\ : std_logic;
signal \N__1292\ : std_logic;
signal \N__1291\ : std_logic;
signal \N__1288\ : std_logic;
signal \N__1283\ : std_logic;
signal \N__1274\ : std_logic;
signal \N__1269\ : std_logic;
signal \N__1266\ : std_logic;
signal \N__1263\ : std_logic;
signal \N__1260\ : std_logic;
signal \N__1257\ : std_logic;
signal \N__1254\ : std_logic;
signal \N__1251\ : std_logic;
signal \N__1248\ : std_logic;
signal \N__1245\ : std_logic;
signal \N__1242\ : std_logic;
signal \N__1239\ : std_logic;
signal \N__1236\ : std_logic;
signal \N__1233\ : std_logic;
signal \N__1230\ : std_logic;
signal \N__1227\ : std_logic;
signal \N__1226\ : std_logic;
signal \N__1225\ : std_logic;
signal \N__1224\ : std_logic;
signal \N__1221\ : std_logic;
signal \N__1218\ : std_logic;
signal \N__1213\ : std_logic;
signal \N__1208\ : std_logic;
signal \N__1203\ : std_logic;
signal \N__1200\ : std_logic;
signal \N__1199\ : std_logic;
signal \N__1198\ : std_logic;
signal \N__1195\ : std_logic;
signal \N__1192\ : std_logic;
signal \N__1189\ : std_logic;
signal \N__1186\ : std_logic;
signal \N__1179\ : std_logic;
signal \N__1176\ : std_logic;
signal \N__1175\ : std_logic;
signal \N__1174\ : std_logic;
signal \N__1171\ : std_logic;
signal \N__1168\ : std_logic;
signal \N__1165\ : std_logic;
signal \N__1158\ : std_logic;
signal \N__1155\ : std_logic;
signal \N__1154\ : std_logic;
signal \N__1151\ : std_logic;
signal \N__1148\ : std_logic;
signal \N__1143\ : std_logic;
signal \N__1140\ : std_logic;
signal \N__1139\ : std_logic;
signal \N__1136\ : std_logic;
signal \N__1133\ : std_logic;
signal \N__1128\ : std_logic;
signal \N__1127\ : std_logic;
signal \N__1122\ : std_logic;
signal \N__1119\ : std_logic;
signal \N__1116\ : std_logic;
signal \N__1113\ : std_logic;
signal \N__1110\ : std_logic;
signal \N__1107\ : std_logic;
signal \N__1104\ : std_logic;
signal \N__1101\ : std_logic;
signal \N__1098\ : std_logic;
signal \N__1095\ : std_logic;
signal \N__1092\ : std_logic;
signal \N__1089\ : std_logic;
signal \N__1086\ : std_logic;
signal \N__1083\ : std_logic;
signal \N__1080\ : std_logic;
signal \N__1077\ : std_logic;
signal \N__1074\ : std_logic;
signal \N__1071\ : std_logic;
signal \N__1068\ : std_logic;
signal \N__1065\ : std_logic;
signal \N__1062\ : std_logic;
signal \N__1059\ : std_logic;
signal \N__1056\ : std_logic;
signal \N__1053\ : std_logic;
signal \N__1050\ : std_logic;
signal \N__1047\ : std_logic;
signal \N__1044\ : std_logic;
signal \N__1041\ : std_logic;
signal \N__1038\ : std_logic;
signal \N__1035\ : std_logic;
signal \N__1032\ : std_logic;
signal \N__1029\ : std_logic;
signal \N__1026\ : std_logic;
signal \N__1023\ : std_logic;
signal \N__1020\ : std_logic;
signal \N__1017\ : std_logic;
signal \N__1014\ : std_logic;
signal \N__1013\ : std_logic;
signal \N__1010\ : std_logic;
signal \N__1009\ : std_logic;
signal \N__1006\ : std_logic;
signal \N__1001\ : std_logic;
signal \N__996\ : std_logic;
signal \N__993\ : std_logic;
signal \N__990\ : std_logic;
signal \N__987\ : std_logic;
signal \N__986\ : std_logic;
signal \N__983\ : std_logic;
signal \N__980\ : std_logic;
signal \N__977\ : std_logic;
signal \N__972\ : std_logic;
signal \N__969\ : std_logic;
signal \N__966\ : std_logic;
signal \N__963\ : std_logic;
signal \N__962\ : std_logic;
signal \N__959\ : std_logic;
signal \N__956\ : std_logic;
signal \N__951\ : std_logic;
signal \N__948\ : std_logic;
signal \N__945\ : std_logic;
signal \N__942\ : std_logic;
signal \N__939\ : std_logic;
signal \N__936\ : std_logic;
signal \N__935\ : std_logic;
signal \N__932\ : std_logic;
signal \N__929\ : std_logic;
signal \N__924\ : std_logic;
signal \N__921\ : std_logic;
signal \N__918\ : std_logic;
signal \N__915\ : std_logic;
signal \N__912\ : std_logic;
signal \N__909\ : std_logic;
signal \N__906\ : std_logic;
signal \N__903\ : std_logic;
signal \N__900\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \oData_c_0\ : std_logic;
signal \oData_c_1\ : std_logic;
signal \pReceive_un12_rstate_3_cascade_\ : std_logic;
signal \N_97_0_i_0_cascade_\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \rCycleCounter_cry_0\ : std_logic;
signal \rCycleCounter_s_2\ : std_logic;
signal \rCycleCounter_cry_1\ : std_logic;
signal \rCycleCounter_s_3\ : std_logic;
signal \rCycleCounter_cry_2\ : std_logic;
signal \rCycleCounterZ0Z_4\ : std_logic;
signal \rCycleCounter_cry_3_THRU_CO\ : std_logic;
signal \rCycleCounter_cry_3\ : std_logic;
signal \rCycleCounterZ0Z_5\ : std_logic;
signal \rCycleCounter_s_5\ : std_logic;
signal \rCycleCounter_cry_4\ : std_logic;
signal \rCycleCounterZ0Z_6\ : std_logic;
signal \rCycleCounter_s_6\ : std_logic;
signal \rCycleCounter_cry_5\ : std_logic;
signal \rCycleCounter_cry_6\ : std_logic;
signal \rCycleCounterZ0Z_7\ : std_logic;
signal \oData_c_5\ : std_logic;
signal \oData_c_2\ : std_logic;
signal \rDatace_1_0_cascade_\ : std_logic;
signal \rData_RNOZ0Z_0\ : std_logic;
signal \rDatace_1_1_cascade_\ : std_logic;
signal \rData_RNOZ0Z_1\ : std_logic;
signal \rDataCounter_0_sqmuxa_cascade_\ : std_logic;
signal \rDataCounter_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \rCycleCounterZ0Z_2\ : std_logic;
signal \rCycleCounterZ0Z_3\ : std_logic;
signal \rCycleCounter_RNIEVAN1Z0Z_0_cascade_\ : std_logic;
signal \pReceive_un12_rstate_4\ : std_logic;
signal \N_97_0_i_cascade_\ : std_logic;
signal \un1_rData_0_sqmuxa_0\ : std_logic;
signal \rDataCounter_0_sqmuxa\ : std_logic;
signal \oData_c_4\ : std_logic;
signal \rDatace_1_4_cascade_\ : std_logic;
signal \rData_RNOZ0Z_4\ : std_logic;
signal \rDatace_1_5_cascade_\ : std_logic;
signal \rData_RNOZ0Z_5\ : std_logic;
signal \rDatace_1_6_cascade_\ : std_logic;
signal \oData_c_6\ : std_logic;
signal \rData_RNOZ0Z_6\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \rDatace_1_2\ : std_logic;
signal \rData_RNOZ0Z_2\ : std_logic;
signal g0_sn : std_logic;
signal \rCycleCounterZ0Z_0\ : std_logic;
signal \N_97_0_i_0\ : std_logic;
signal \rCycleCounter_cry_0_THRU_CO\ : std_logic;
signal \rCycleCounterZ0Z_1\ : std_logic;
signal \pReceive_rstate\ : std_logic;
signal \CO0_0\ : std_logic;
signal \rCycleCountere_0_i\ : std_logic;
signal \rState_0_repZ0Z1\ : std_logic;
signal \rDataCounterZ0Z_2\ : std_logic;
signal \rDataCounterZ0Z_1\ : std_logic;
signal \rDataCounterZ0Z_0\ : std_logic;
signal \rState_1_repZ0Z1\ : std_logic;
signal \rDatace_0_3_cascade_\ : std_logic;
signal \oData_c_3\ : std_logic;
signal \rData_RNOZ0Z_3\ : std_logic;
signal \oDataReady_c\ : std_logic;
signal \pReceive_rdata_7\ : std_logic;
signal \N_97_0_i\ : std_logic;
signal \rStateZ0Z_0\ : std_logic;
signal \rState_fastZ0Z_1\ : std_logic;
signal \rStateZ0Z_1\ : std_logic;
signal \rState_fastZ0Z_0\ : std_logic;
signal \un1_rCycleCounter_2_sqmuxa_0\ : std_logic;
signal \iSerial_c\ : std_logic;
signal \oData_c_7\ : std_logic;
signal \iClk_c_g\ : std_logic;
signal \rData_RNOZ0Z_7\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \iClk_wire\ : std_logic;
signal \oData_wire\ : std_logic_vector(7 downto 0);
signal \oDataReady_wire\ : std_logic;
signal \iSerial_wire\ : std_logic;

begin
    \iClk_wire\ <= iClk;
    oData <= \oData_wire\;
    oDataReady <= \oDataReady_wire\;
    \iSerial_wire\ <= iSerial;

    \iClk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2410\,
            GLOBALBUFFEROUTPUT => \iClk_c_g\
        );

    \iClk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2412\,
            DIN => \N__2411\,
            DOUT => \N__2410\,
            PACKAGEPIN => \iClk_wire\
        );

    \iClk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2412\,
            PADOUT => \N__2411\,
            PADIN => \N__2410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oData_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2401\,
            DIN => \N__2400\,
            DOUT => \N__2399\,
            PACKAGEPIN => \oData_wire\(3)
        );

    \oData_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2401\,
            PADOUT => \N__2400\,
            PADIN => \N__2399\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2301\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oDataReady_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2392\,
            DIN => \N__2391\,
            DOUT => \N__2390\,
            PACKAGEPIN => \oDataReady_wire\
        );

    \oDataReady_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2392\,
            PADOUT => \N__2391\,
            PADIN => \N__2390\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2283\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oData_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2383\,
            DIN => \N__2382\,
            DOUT => \N__2381\,
            PACKAGEPIN => \oData_wire\(4)
        );

    \oData_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2383\,
            PADOUT => \N__2382\,
            PADIN => \N__2381\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1119\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oData_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2374\,
            DIN => \N__2373\,
            DOUT => \N__2372\,
            PACKAGEPIN => \oData_wire\(2)
        );

    \oData_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2374\,
            PADOUT => \N__2373\,
            PADIN => \N__2372\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1074\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oData_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2365\,
            DIN => \N__2364\,
            DOUT => \N__2363\,
            PACKAGEPIN => \oData_wire\(0)
        );

    \oData_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2365\,
            PADOUT => \N__2364\,
            PADIN => \N__2363\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__903\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iSerial_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2356\,
            DIN => \N__2355\,
            DOUT => \N__2354\,
            PACKAGEPIN => \iSerial_wire\
        );

    \iSerial_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2356\,
            PADOUT => \N__2355\,
            PADIN => \N__2354\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iSerial_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oData_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2347\,
            DIN => \N__2346\,
            DOUT => \N__2345\,
            PACKAGEPIN => \oData_wire\(7)
        );

    \oData_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2347\,
            PADOUT => \N__2346\,
            PADIN => \N__2345\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1842\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oData_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2338\,
            DIN => \N__2337\,
            DOUT => \N__2336\,
            PACKAGEPIN => \oData_wire\(5)
        );

    \oData_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2338\,
            PADOUT => \N__2337\,
            PADIN => \N__2336\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__924\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oData_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2329\,
            DIN => \N__2328\,
            DOUT => \N__2327\,
            PACKAGEPIN => \oData_wire\(1)
        );

    \oData_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2329\,
            PADOUT => \N__2328\,
            PADIN => \N__2327\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__915\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oData_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2320\,
            DIN => \N__2319\,
            DOUT => \N__2318\,
            PACKAGEPIN => \oData_wire\(6)
        );

    \oData_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2320\,
            PADOUT => \N__2319\,
            PADIN => \N__2318\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1329\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__545\ : IoInMux
    port map (
            O => \N__2301\,
            I => \N__2298\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__2298\,
            I => \N__2295\
        );

    \I__543\ : Odrv12
    port map (
            O => \N__2295\,
            I => \oData_c_3\
        );

    \I__542\ : CEMux
    port map (
            O => \N__2292\,
            I => \N__2289\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__2289\,
            I => \N__2286\
        );

    \I__540\ : Odrv4
    port map (
            O => \N__2286\,
            I => \rData_RNOZ0Z_3\
        );

    \I__539\ : IoInMux
    port map (
            O => \N__2283\,
            I => \N__2280\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__2280\,
            I => \N__2277\
        );

    \I__537\ : IoSpan4Mux
    port map (
            O => \N__2277\,
            I => \N__2274\
        );

    \I__536\ : Span4Mux_s3_h
    port map (
            O => \N__2274\,
            I => \N__2270\
        );

    \I__535\ : InMux
    port map (
            O => \N__2273\,
            I => \N__2267\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__2270\,
            I => \oDataReady_c\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2267\,
            I => \oDataReady_c\
        );

    \I__532\ : InMux
    port map (
            O => \N__2262\,
            I => \N__2256\
        );

    \I__531\ : InMux
    port map (
            O => \N__2261\,
            I => \N__2256\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__2256\,
            I => \N__2253\
        );

    \I__529\ : Span4Mux_h
    port map (
            O => \N__2253\,
            I => \N__2249\
        );

    \I__528\ : InMux
    port map (
            O => \N__2252\,
            I => \N__2246\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__2249\,
            I => \pReceive_rdata_7\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__2246\,
            I => \pReceive_rdata_7\
        );

    \I__525\ : InMux
    port map (
            O => \N__2241\,
            I => \N__2236\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__2240\,
            I => \N__2233\
        );

    \I__523\ : InMux
    port map (
            O => \N__2239\,
            I => \N__2220\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__2236\,
            I => \N__2217\
        );

    \I__521\ : InMux
    port map (
            O => \N__2233\,
            I => \N__2212\
        );

    \I__520\ : InMux
    port map (
            O => \N__2232\,
            I => \N__2212\
        );

    \I__519\ : InMux
    port map (
            O => \N__2231\,
            I => \N__2203\
        );

    \I__518\ : InMux
    port map (
            O => \N__2230\,
            I => \N__2203\
        );

    \I__517\ : InMux
    port map (
            O => \N__2229\,
            I => \N__2203\
        );

    \I__516\ : InMux
    port map (
            O => \N__2228\,
            I => \N__2203\
        );

    \I__515\ : InMux
    port map (
            O => \N__2227\,
            I => \N__2198\
        );

    \I__514\ : InMux
    port map (
            O => \N__2226\,
            I => \N__2198\
        );

    \I__513\ : InMux
    port map (
            O => \N__2225\,
            I => \N__2191\
        );

    \I__512\ : InMux
    port map (
            O => \N__2224\,
            I => \N__2191\
        );

    \I__511\ : InMux
    port map (
            O => \N__2223\,
            I => \N__2191\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__2220\,
            I => \N__2188\
        );

    \I__509\ : Span4Mux_h
    port map (
            O => \N__2217\,
            I => \N__2185\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__2212\,
            I => \N__2182\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__2203\,
            I => \N_97_0_i\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__2198\,
            I => \N_97_0_i\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__2191\,
            I => \N_97_0_i\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__2188\,
            I => \N_97_0_i\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__2185\,
            I => \N_97_0_i\
        );

    \I__502\ : Odrv12
    port map (
            O => \N__2182\,
            I => \N_97_0_i\
        );

    \I__501\ : InMux
    port map (
            O => \N__2169\,
            I => \N__2164\
        );

    \I__500\ : InMux
    port map (
            O => \N__2168\,
            I => \N__2158\
        );

    \I__499\ : InMux
    port map (
            O => \N__2167\,
            I => \N__2155\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__2164\,
            I => \N__2147\
        );

    \I__497\ : InMux
    port map (
            O => \N__2163\,
            I => \N__2140\
        );

    \I__496\ : InMux
    port map (
            O => \N__2162\,
            I => \N__2140\
        );

    \I__495\ : InMux
    port map (
            O => \N__2161\,
            I => \N__2140\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2158\,
            I => \N__2134\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__2155\,
            I => \N__2134\
        );

    \I__492\ : InMux
    port map (
            O => \N__2154\,
            I => \N__2129\
        );

    \I__491\ : InMux
    port map (
            O => \N__2153\,
            I => \N__2129\
        );

    \I__490\ : InMux
    port map (
            O => \N__2152\,
            I => \N__2122\
        );

    \I__489\ : InMux
    port map (
            O => \N__2151\,
            I => \N__2122\
        );

    \I__488\ : InMux
    port map (
            O => \N__2150\,
            I => \N__2122\
        );

    \I__487\ : Span4Mux_v
    port map (
            O => \N__2147\,
            I => \N__2117\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__2140\,
            I => \N__2117\
        );

    \I__485\ : InMux
    port map (
            O => \N__2139\,
            I => \N__2114\
        );

    \I__484\ : Odrv4
    port map (
            O => \N__2134\,
            I => \rStateZ0Z_0\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2129\,
            I => \rStateZ0Z_0\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__2122\,
            I => \rStateZ0Z_0\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__2117\,
            I => \rStateZ0Z_0\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2114\,
            I => \rStateZ0Z_0\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__2103\,
            I => \N__2098\
        );

    \I__478\ : InMux
    port map (
            O => \N__2102\,
            I => \N__2095\
        );

    \I__477\ : InMux
    port map (
            O => \N__2101\,
            I => \N__2090\
        );

    \I__476\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2090\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2095\,
            I => \rState_fastZ0Z_1\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2090\,
            I => \rState_fastZ0Z_1\
        );

    \I__473\ : InMux
    port map (
            O => \N__2085\,
            I => \N__2079\
        );

    \I__472\ : InMux
    port map (
            O => \N__2084\,
            I => \N__2079\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__2079\,
            I => \N__2074\
        );

    \I__470\ : InMux
    port map (
            O => \N__2078\,
            I => \N__2069\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__2077\,
            I => \N__2061\
        );

    \I__468\ : Span4Mux_v
    port map (
            O => \N__2074\,
            I => \N__2058\
        );

    \I__467\ : InMux
    port map (
            O => \N__2073\,
            I => \N__2053\
        );

    \I__466\ : InMux
    port map (
            O => \N__2072\,
            I => \N__2053\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__2069\,
            I => \N__2050\
        );

    \I__464\ : InMux
    port map (
            O => \N__2068\,
            I => \N__2043\
        );

    \I__463\ : InMux
    port map (
            O => \N__2067\,
            I => \N__2043\
        );

    \I__462\ : InMux
    port map (
            O => \N__2066\,
            I => \N__2043\
        );

    \I__461\ : InMux
    port map (
            O => \N__2065\,
            I => \N__2036\
        );

    \I__460\ : InMux
    port map (
            O => \N__2064\,
            I => \N__2036\
        );

    \I__459\ : InMux
    port map (
            O => \N__2061\,
            I => \N__2036\
        );

    \I__458\ : Span4Mux_s0_h
    port map (
            O => \N__2058\,
            I => \N__2031\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2053\,
            I => \N__2031\
        );

    \I__456\ : Odrv4
    port map (
            O => \N__2050\,
            I => \rStateZ0Z_1\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2043\,
            I => \rStateZ0Z_1\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2036\,
            I => \rStateZ0Z_1\
        );

    \I__453\ : Odrv4
    port map (
            O => \N__2031\,
            I => \rStateZ0Z_1\
        );

    \I__452\ : InMux
    port map (
            O => \N__2022\,
            I => \N__2017\
        );

    \I__451\ : InMux
    port map (
            O => \N__2021\,
            I => \N__2012\
        );

    \I__450\ : InMux
    port map (
            O => \N__2020\,
            I => \N__2012\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2017\,
            I => \rState_fastZ0Z_0\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2012\,
            I => \rState_fastZ0Z_0\
        );

    \I__447\ : CEMux
    port map (
            O => \N__2007\,
            I => \N__2002\
        );

    \I__446\ : CEMux
    port map (
            O => \N__2006\,
            I => \N__1999\
        );

    \I__445\ : CEMux
    port map (
            O => \N__2005\,
            I => \N__1996\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2002\,
            I => \un1_rCycleCounter_2_sqmuxa_0\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__1999\,
            I => \un1_rCycleCounter_2_sqmuxa_0\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__1996\,
            I => \un1_rCycleCounter_2_sqmuxa_0\
        );

    \I__441\ : CascadeMux
    port map (
            O => \N__1989\,
            I => \N__1983\
        );

    \I__440\ : InMux
    port map (
            O => \N__1988\,
            I => \N__1979\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__1987\,
            I => \N__1975\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__1986\,
            I => \N__1971\
        );

    \I__437\ : InMux
    port map (
            O => \N__1983\,
            I => \N__1961\
        );

    \I__436\ : InMux
    port map (
            O => \N__1982\,
            I => \N__1961\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__1979\,
            I => \N__1958\
        );

    \I__434\ : InMux
    port map (
            O => \N__1978\,
            I => \N__1955\
        );

    \I__433\ : InMux
    port map (
            O => \N__1975\,
            I => \N__1948\
        );

    \I__432\ : InMux
    port map (
            O => \N__1974\,
            I => \N__1948\
        );

    \I__431\ : InMux
    port map (
            O => \N__1971\,
            I => \N__1948\
        );

    \I__430\ : InMux
    port map (
            O => \N__1970\,
            I => \N__1945\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__1969\,
            I => \N__1941\
        );

    \I__428\ : CascadeMux
    port map (
            O => \N__1968\,
            I => \N__1938\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__1967\,
            I => \N__1935\
        );

    \I__426\ : InMux
    port map (
            O => \N__1966\,
            I => \N__1929\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__1961\,
            I => \N__1924\
        );

    \I__424\ : Span4Mux_v
    port map (
            O => \N__1958\,
            I => \N__1915\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__1955\,
            I => \N__1915\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__1948\,
            I => \N__1915\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__1945\,
            I => \N__1915\
        );

    \I__420\ : InMux
    port map (
            O => \N__1944\,
            I => \N__1912\
        );

    \I__419\ : InMux
    port map (
            O => \N__1941\,
            I => \N__1905\
        );

    \I__418\ : InMux
    port map (
            O => \N__1938\,
            I => \N__1905\
        );

    \I__417\ : InMux
    port map (
            O => \N__1935\,
            I => \N__1905\
        );

    \I__416\ : InMux
    port map (
            O => \N__1934\,
            I => \N__1902\
        );

    \I__415\ : InMux
    port map (
            O => \N__1933\,
            I => \N__1899\
        );

    \I__414\ : InMux
    port map (
            O => \N__1932\,
            I => \N__1895\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__1929\,
            I => \N__1892\
        );

    \I__412\ : InMux
    port map (
            O => \N__1928\,
            I => \N__1889\
        );

    \I__411\ : InMux
    port map (
            O => \N__1927\,
            I => \N__1886\
        );

    \I__410\ : Span4Mux_v
    port map (
            O => \N__1924\,
            I => \N__1881\
        );

    \I__409\ : Span4Mux_v
    port map (
            O => \N__1915\,
            I => \N__1881\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__1912\,
            I => \N__1872\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__1905\,
            I => \N__1872\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__1902\,
            I => \N__1872\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__1899\,
            I => \N__1872\
        );

    \I__404\ : InMux
    port map (
            O => \N__1898\,
            I => \N__1869\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__1895\,
            I => \N__1860\
        );

    \I__402\ : Sp12to4
    port map (
            O => \N__1892\,
            I => \N__1860\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__1889\,
            I => \N__1860\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__1886\,
            I => \N__1860\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__1881\,
            I => \N__1853\
        );

    \I__398\ : Span4Mux_v
    port map (
            O => \N__1872\,
            I => \N__1853\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__1869\,
            I => \N__1853\
        );

    \I__396\ : Span12Mux_v
    port map (
            O => \N__1860\,
            I => \N__1850\
        );

    \I__395\ : Span4Mux_v
    port map (
            O => \N__1853\,
            I => \N__1847\
        );

    \I__394\ : Odrv12
    port map (
            O => \N__1850\,
            I => \iSerial_c\
        );

    \I__393\ : Odrv4
    port map (
            O => \N__1847\,
            I => \iSerial_c\
        );

    \I__392\ : IoInMux
    port map (
            O => \N__1842\,
            I => \N__1839\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__1839\,
            I => \N__1836\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__1836\,
            I => \oData_c_7\
        );

    \I__389\ : ClkMux
    port map (
            O => \N__1833\,
            I => \N__1785\
        );

    \I__388\ : ClkMux
    port map (
            O => \N__1832\,
            I => \N__1785\
        );

    \I__387\ : ClkMux
    port map (
            O => \N__1831\,
            I => \N__1785\
        );

    \I__386\ : ClkMux
    port map (
            O => \N__1830\,
            I => \N__1785\
        );

    \I__385\ : ClkMux
    port map (
            O => \N__1829\,
            I => \N__1785\
        );

    \I__384\ : ClkMux
    port map (
            O => \N__1828\,
            I => \N__1785\
        );

    \I__383\ : ClkMux
    port map (
            O => \N__1827\,
            I => \N__1785\
        );

    \I__382\ : ClkMux
    port map (
            O => \N__1826\,
            I => \N__1785\
        );

    \I__381\ : ClkMux
    port map (
            O => \N__1825\,
            I => \N__1785\
        );

    \I__380\ : ClkMux
    port map (
            O => \N__1824\,
            I => \N__1785\
        );

    \I__379\ : ClkMux
    port map (
            O => \N__1823\,
            I => \N__1785\
        );

    \I__378\ : ClkMux
    port map (
            O => \N__1822\,
            I => \N__1785\
        );

    \I__377\ : ClkMux
    port map (
            O => \N__1821\,
            I => \N__1785\
        );

    \I__376\ : ClkMux
    port map (
            O => \N__1820\,
            I => \N__1785\
        );

    \I__375\ : ClkMux
    port map (
            O => \N__1819\,
            I => \N__1785\
        );

    \I__374\ : ClkMux
    port map (
            O => \N__1818\,
            I => \N__1785\
        );

    \I__373\ : GlobalMux
    port map (
            O => \N__1785\,
            I => \N__1782\
        );

    \I__372\ : gio2CtrlBuf
    port map (
            O => \N__1782\,
            I => \iClk_c_g\
        );

    \I__371\ : CEMux
    port map (
            O => \N__1779\,
            I => \N__1776\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__1776\,
            I => \N__1773\
        );

    \I__369\ : Span4Mux_v
    port map (
            O => \N__1773\,
            I => \N__1770\
        );

    \I__368\ : Odrv4
    port map (
            O => \N__1770\,
            I => \rData_RNOZ0Z_7\
        );

    \I__367\ : InMux
    port map (
            O => \N__1767\,
            I => \N__1761\
        );

    \I__366\ : InMux
    port map (
            O => \N__1766\,
            I => \N__1761\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__1761\,
            I => \N__1753\
        );

    \I__364\ : InMux
    port map (
            O => \N__1760\,
            I => \N__1750\
        );

    \I__363\ : InMux
    port map (
            O => \N__1759\,
            I => \N__1741\
        );

    \I__362\ : InMux
    port map (
            O => \N__1758\,
            I => \N__1741\
        );

    \I__361\ : InMux
    port map (
            O => \N__1757\,
            I => \N__1741\
        );

    \I__360\ : InMux
    port map (
            O => \N__1756\,
            I => \N__1741\
        );

    \I__359\ : Odrv4
    port map (
            O => \N__1753\,
            I => \N_97_0_i_0\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__1750\,
            I => \N_97_0_i_0\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__1741\,
            I => \N_97_0_i_0\
        );

    \I__356\ : InMux
    port map (
            O => \N__1734\,
            I => \N__1731\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__1731\,
            I => \N__1728\
        );

    \I__354\ : Span4Mux_v
    port map (
            O => \N__1728\,
            I => \N__1725\
        );

    \I__353\ : Odrv4
    port map (
            O => \N__1725\,
            I => \rCycleCounter_cry_0_THRU_CO\
        );

    \I__352\ : InMux
    port map (
            O => \N__1722\,
            I => \N__1719\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__1719\,
            I => \N__1713\
        );

    \I__350\ : InMux
    port map (
            O => \N__1718\,
            I => \N__1710\
        );

    \I__349\ : InMux
    port map (
            O => \N__1717\,
            I => \N__1705\
        );

    \I__348\ : InMux
    port map (
            O => \N__1716\,
            I => \N__1705\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__1713\,
            I => \N__1700\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__1710\,
            I => \N__1700\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__1705\,
            I => \rCycleCounterZ0Z_1\
        );

    \I__344\ : Odrv4
    port map (
            O => \N__1700\,
            I => \rCycleCounterZ0Z_1\
        );

    \I__343\ : SRMux
    port map (
            O => \N__1695\,
            I => \N__1692\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__1692\,
            I => \N__1686\
        );

    \I__341\ : InMux
    port map (
            O => \N__1691\,
            I => \N__1679\
        );

    \I__340\ : InMux
    port map (
            O => \N__1690\,
            I => \N__1679\
        );

    \I__339\ : InMux
    port map (
            O => \N__1689\,
            I => \N__1679\
        );

    \I__338\ : Span4Mux_h
    port map (
            O => \N__1686\,
            I => \N__1676\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__1679\,
            I => \N__1673\
        );

    \I__336\ : Odrv4
    port map (
            O => \N__1676\,
            I => \pReceive_rstate\
        );

    \I__335\ : Odrv4
    port map (
            O => \N__1673\,
            I => \pReceive_rstate\
        );

    \I__334\ : InMux
    port map (
            O => \N__1668\,
            I => \N__1664\
        );

    \I__333\ : InMux
    port map (
            O => \N__1667\,
            I => \N__1661\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__1664\,
            I => \N__1656\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__1661\,
            I => \N__1656\
        );

    \I__330\ : Odrv4
    port map (
            O => \N__1656\,
            I => \CO0_0\
        );

    \I__329\ : CEMux
    port map (
            O => \N__1653\,
            I => \N__1649\
        );

    \I__328\ : CEMux
    port map (
            O => \N__1652\,
            I => \N__1646\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__1649\,
            I => \N__1643\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__1646\,
            I => \N__1640\
        );

    \I__325\ : Span4Mux_v
    port map (
            O => \N__1643\,
            I => \N__1635\
        );

    \I__324\ : Span4Mux_s1_h
    port map (
            O => \N__1640\,
            I => \N__1635\
        );

    \I__323\ : Span4Mux_h
    port map (
            O => \N__1635\,
            I => \N__1631\
        );

    \I__322\ : CEMux
    port map (
            O => \N__1634\,
            I => \N__1628\
        );

    \I__321\ : Span4Mux_s1_h
    port map (
            O => \N__1631\,
            I => \N__1623\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__1628\,
            I => \N__1623\
        );

    \I__319\ : Odrv4
    port map (
            O => \N__1623\,
            I => \rCycleCountere_0_i\
        );

    \I__318\ : InMux
    port map (
            O => \N__1620\,
            I => \N__1614\
        );

    \I__317\ : InMux
    port map (
            O => \N__1619\,
            I => \N__1614\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1614\,
            I => \N__1608\
        );

    \I__315\ : InMux
    port map (
            O => \N__1613\,
            I => \N__1605\
        );

    \I__314\ : InMux
    port map (
            O => \N__1612\,
            I => \N__1600\
        );

    \I__313\ : InMux
    port map (
            O => \N__1611\,
            I => \N__1600\
        );

    \I__312\ : Span4Mux_v
    port map (
            O => \N__1608\,
            I => \N__1596\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__1605\,
            I => \N__1591\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__1600\,
            I => \N__1588\
        );

    \I__309\ : InMux
    port map (
            O => \N__1599\,
            I => \N__1585\
        );

    \I__308\ : Span4Mux_s1_h
    port map (
            O => \N__1596\,
            I => \N__1582\
        );

    \I__307\ : InMux
    port map (
            O => \N__1595\,
            I => \N__1577\
        );

    \I__306\ : InMux
    port map (
            O => \N__1594\,
            I => \N__1577\
        );

    \I__305\ : Span4Mux_s3_h
    port map (
            O => \N__1591\,
            I => \N__1572\
        );

    \I__304\ : Span4Mux_s3_h
    port map (
            O => \N__1588\,
            I => \N__1572\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__1585\,
            I => \rState_0_repZ0Z1\
        );

    \I__302\ : Odrv4
    port map (
            O => \N__1582\,
            I => \rState_0_repZ0Z1\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__1577\,
            I => \rState_0_repZ0Z1\
        );

    \I__300\ : Odrv4
    port map (
            O => \N__1572\,
            I => \rState_0_repZ0Z1\
        );

    \I__299\ : InMux
    port map (
            O => \N__1563\,
            I => \N__1559\
        );

    \I__298\ : CascadeMux
    port map (
            O => \N__1562\,
            I => \N__1553\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__1559\,
            I => \N__1550\
        );

    \I__296\ : InMux
    port map (
            O => \N__1558\,
            I => \N__1543\
        );

    \I__295\ : InMux
    port map (
            O => \N__1557\,
            I => \N__1543\
        );

    \I__294\ : InMux
    port map (
            O => \N__1556\,
            I => \N__1543\
        );

    \I__293\ : InMux
    port map (
            O => \N__1553\,
            I => \N__1536\
        );

    \I__292\ : Span4Mux_v
    port map (
            O => \N__1550\,
            I => \N__1533\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1543\,
            I => \N__1530\
        );

    \I__290\ : InMux
    port map (
            O => \N__1542\,
            I => \N__1521\
        );

    \I__289\ : InMux
    port map (
            O => \N__1541\,
            I => \N__1521\
        );

    \I__288\ : InMux
    port map (
            O => \N__1540\,
            I => \N__1521\
        );

    \I__287\ : InMux
    port map (
            O => \N__1539\,
            I => \N__1521\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1536\,
            I => \rDataCounterZ0Z_2\
        );

    \I__285\ : Odrv4
    port map (
            O => \N__1533\,
            I => \rDataCounterZ0Z_2\
        );

    \I__284\ : Odrv4
    port map (
            O => \N__1530\,
            I => \rDataCounterZ0Z_2\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__1521\,
            I => \rDataCounterZ0Z_2\
        );

    \I__282\ : InMux
    port map (
            O => \N__1512\,
            I => \N__1509\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__1509\,
            I => \N__1504\
        );

    \I__280\ : InMux
    port map (
            O => \N__1508\,
            I => \N__1492\
        );

    \I__279\ : InMux
    port map (
            O => \N__1507\,
            I => \N__1492\
        );

    \I__278\ : Span4Mux_h
    port map (
            O => \N__1504\,
            I => \N__1489\
        );

    \I__277\ : InMux
    port map (
            O => \N__1503\,
            I => \N__1482\
        );

    \I__276\ : InMux
    port map (
            O => \N__1502\,
            I => \N__1482\
        );

    \I__275\ : InMux
    port map (
            O => \N__1501\,
            I => \N__1482\
        );

    \I__274\ : InMux
    port map (
            O => \N__1500\,
            I => \N__1473\
        );

    \I__273\ : InMux
    port map (
            O => \N__1499\,
            I => \N__1473\
        );

    \I__272\ : InMux
    port map (
            O => \N__1498\,
            I => \N__1473\
        );

    \I__271\ : InMux
    port map (
            O => \N__1497\,
            I => \N__1473\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__1492\,
            I => \rDataCounterZ0Z_1\
        );

    \I__269\ : Odrv4
    port map (
            O => \N__1489\,
            I => \rDataCounterZ0Z_1\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1482\,
            I => \rDataCounterZ0Z_1\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__1473\,
            I => \rDataCounterZ0Z_1\
        );

    \I__266\ : InMux
    port map (
            O => \N__1464\,
            I => \N__1459\
        );

    \I__265\ : CascadeMux
    port map (
            O => \N__1463\,
            I => \N__1456\
        );

    \I__264\ : InMux
    port map (
            O => \N__1462\,
            I => \N__1453\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1459\,
            I => \N__1450\
        );

    \I__262\ : InMux
    port map (
            O => \N__1456\,
            I => \N__1440\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__1453\,
            I => \N__1437\
        );

    \I__260\ : Span4Mux_h
    port map (
            O => \N__1450\,
            I => \N__1434\
        );

    \I__259\ : InMux
    port map (
            O => \N__1449\,
            I => \N__1427\
        );

    \I__258\ : InMux
    port map (
            O => \N__1448\,
            I => \N__1427\
        );

    \I__257\ : InMux
    port map (
            O => \N__1447\,
            I => \N__1427\
        );

    \I__256\ : InMux
    port map (
            O => \N__1446\,
            I => \N__1418\
        );

    \I__255\ : InMux
    port map (
            O => \N__1445\,
            I => \N__1418\
        );

    \I__254\ : InMux
    port map (
            O => \N__1444\,
            I => \N__1418\
        );

    \I__253\ : InMux
    port map (
            O => \N__1443\,
            I => \N__1418\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__1440\,
            I => \rDataCounterZ0Z_0\
        );

    \I__251\ : Odrv12
    port map (
            O => \N__1437\,
            I => \rDataCounterZ0Z_0\
        );

    \I__250\ : Odrv4
    port map (
            O => \N__1434\,
            I => \rDataCounterZ0Z_0\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1427\,
            I => \rDataCounterZ0Z_0\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1418\,
            I => \rDataCounterZ0Z_0\
        );

    \I__247\ : CascadeMux
    port map (
            O => \N__1407\,
            I => \N__1403\
        );

    \I__246\ : CascadeMux
    port map (
            O => \N__1406\,
            I => \N__1399\
        );

    \I__245\ : InMux
    port map (
            O => \N__1403\,
            I => \N__1394\
        );

    \I__244\ : InMux
    port map (
            O => \N__1402\,
            I => \N__1391\
        );

    \I__243\ : InMux
    port map (
            O => \N__1399\,
            I => \N__1386\
        );

    \I__242\ : InMux
    port map (
            O => \N__1398\,
            I => \N__1383\
        );

    \I__241\ : InMux
    port map (
            O => \N__1397\,
            I => \N__1379\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__1394\,
            I => \N__1374\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1391\,
            I => \N__1374\
        );

    \I__238\ : InMux
    port map (
            O => \N__1390\,
            I => \N__1369\
        );

    \I__237\ : InMux
    port map (
            O => \N__1389\,
            I => \N__1369\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__1386\,
            I => \N__1363\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1383\,
            I => \N__1363\
        );

    \I__234\ : InMux
    port map (
            O => \N__1382\,
            I => \N__1360\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1379\,
            I => \N__1357\
        );

    \I__232\ : Span4Mux_v
    port map (
            O => \N__1374\,
            I => \N__1352\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1369\,
            I => \N__1352\
        );

    \I__230\ : InMux
    port map (
            O => \N__1368\,
            I => \N__1349\
        );

    \I__229\ : Span4Mux_s3_h
    port map (
            O => \N__1363\,
            I => \N__1346\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1360\,
            I => \rState_1_repZ0Z1\
        );

    \I__227\ : Odrv4
    port map (
            O => \N__1357\,
            I => \rState_1_repZ0Z1\
        );

    \I__226\ : Odrv4
    port map (
            O => \N__1352\,
            I => \rState_1_repZ0Z1\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__1349\,
            I => \rState_1_repZ0Z1\
        );

    \I__224\ : Odrv4
    port map (
            O => \N__1346\,
            I => \rState_1_repZ0Z1\
        );

    \I__223\ : CascadeMux
    port map (
            O => \N__1335\,
            I => \rDatace_0_3_cascade_\
        );

    \I__222\ : CascadeMux
    port map (
            O => \N__1332\,
            I => \rDatace_1_6_cascade_\
        );

    \I__221\ : IoInMux
    port map (
            O => \N__1329\,
            I => \N__1326\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__1326\,
            I => \N__1323\
        );

    \I__219\ : Span4Mux_s1_v
    port map (
            O => \N__1323\,
            I => \N__1320\
        );

    \I__218\ : Odrv4
    port map (
            O => \N__1320\,
            I => \oData_c_6\
        );

    \I__217\ : CEMux
    port map (
            O => \N__1317\,
            I => \N__1314\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__1314\,
            I => \N__1311\
        );

    \I__215\ : Odrv12
    port map (
            O => \N__1311\,
            I => \rData_RNOZ0Z_6\
        );

    \I__214\ : CascadeMux
    port map (
            O => \N__1308\,
            I => \N__1301\
        );

    \I__213\ : CascadeMux
    port map (
            O => \N__1307\,
            I => \N__1298\
        );

    \I__212\ : CascadeMux
    port map (
            O => \N__1306\,
            I => \N__1295\
        );

    \I__211\ : CascadeMux
    port map (
            O => \N__1305\,
            I => \N__1292\
        );

    \I__210\ : CascadeMux
    port map (
            O => \N__1304\,
            I => \N__1288\
        );

    \I__209\ : InMux
    port map (
            O => \N__1301\,
            I => \N__1283\
        );

    \I__208\ : InMux
    port map (
            O => \N__1298\,
            I => \N__1283\
        );

    \I__207\ : InMux
    port map (
            O => \N__1295\,
            I => \N__1274\
        );

    \I__206\ : InMux
    port map (
            O => \N__1292\,
            I => \N__1274\
        );

    \I__205\ : InMux
    port map (
            O => \N__1291\,
            I => \N__1274\
        );

    \I__204\ : InMux
    port map (
            O => \N__1288\,
            I => \N__1274\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__1283\,
            I => \N__1269\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1274\,
            I => \N__1269\
        );

    \I__201\ : Span4Mux_v
    port map (
            O => \N__1269\,
            I => \N__1266\
        );

    \I__200\ : Odrv4
    port map (
            O => \N__1266\,
            I => \CONSTANT_ONE_NET\
        );

    \I__199\ : InMux
    port map (
            O => \N__1263\,
            I => \N__1260\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1260\,
            I => \N__1257\
        );

    \I__197\ : Odrv12
    port map (
            O => \N__1257\,
            I => \rDatace_1_2\
        );

    \I__196\ : CEMux
    port map (
            O => \N__1254\,
            I => \N__1251\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1251\,
            I => \N__1248\
        );

    \I__194\ : Span4Mux_s2_h
    port map (
            O => \N__1248\,
            I => \N__1245\
        );

    \I__193\ : Odrv4
    port map (
            O => \N__1245\,
            I => \rData_RNOZ0Z_2\
        );

    \I__192\ : InMux
    port map (
            O => \N__1242\,
            I => \N__1239\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1239\,
            I => \N__1236\
        );

    \I__190\ : Odrv12
    port map (
            O => \N__1236\,
            I => g0_sn
        );

    \I__189\ : CascadeMux
    port map (
            O => \N__1233\,
            I => \N__1230\
        );

    \I__188\ : InMux
    port map (
            O => \N__1230\,
            I => \N__1227\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1227\,
            I => \N__1221\
        );

    \I__186\ : InMux
    port map (
            O => \N__1226\,
            I => \N__1218\
        );

    \I__185\ : InMux
    port map (
            O => \N__1225\,
            I => \N__1213\
        );

    \I__184\ : InMux
    port map (
            O => \N__1224\,
            I => \N__1213\
        );

    \I__183\ : Span4Mux_v
    port map (
            O => \N__1221\,
            I => \N__1208\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__1218\,
            I => \N__1208\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1213\,
            I => \rCycleCounterZ0Z_0\
        );

    \I__180\ : Odrv4
    port map (
            O => \N__1208\,
            I => \rCycleCounterZ0Z_0\
        );

    \I__179\ : CascadeMux
    port map (
            O => \N__1203\,
            I => \N__1200\
        );

    \I__178\ : InMux
    port map (
            O => \N__1200\,
            I => \N__1195\
        );

    \I__177\ : InMux
    port map (
            O => \N__1199\,
            I => \N__1192\
        );

    \I__176\ : InMux
    port map (
            O => \N__1198\,
            I => \N__1189\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1195\,
            I => \N__1186\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1192\,
            I => \rCycleCounterZ0Z_2\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1189\,
            I => \rCycleCounterZ0Z_2\
        );

    \I__172\ : Odrv4
    port map (
            O => \N__1186\,
            I => \rCycleCounterZ0Z_2\
        );

    \I__171\ : CascadeMux
    port map (
            O => \N__1179\,
            I => \N__1176\
        );

    \I__170\ : InMux
    port map (
            O => \N__1176\,
            I => \N__1171\
        );

    \I__169\ : InMux
    port map (
            O => \N__1175\,
            I => \N__1168\
        );

    \I__168\ : InMux
    port map (
            O => \N__1174\,
            I => \N__1165\
        );

    \I__167\ : LocalMux
    port map (
            O => \N__1171\,
            I => \rCycleCounterZ0Z_3\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1168\,
            I => \rCycleCounterZ0Z_3\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__1165\,
            I => \rCycleCounterZ0Z_3\
        );

    \I__164\ : CascadeMux
    port map (
            O => \N__1158\,
            I => \rCycleCounter_RNIEVAN1Z0Z_0_cascade_\
        );

    \I__163\ : InMux
    port map (
            O => \N__1155\,
            I => \N__1151\
        );

    \I__162\ : InMux
    port map (
            O => \N__1154\,
            I => \N__1148\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1151\,
            I => \pReceive_un12_rstate_4\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1148\,
            I => \pReceive_un12_rstate_4\
        );

    \I__159\ : CascadeMux
    port map (
            O => \N__1143\,
            I => \N_97_0_i_cascade_\
        );

    \I__158\ : InMux
    port map (
            O => \N__1140\,
            I => \N__1136\
        );

    \I__157\ : InMux
    port map (
            O => \N__1139\,
            I => \N__1133\
        );

    \I__156\ : LocalMux
    port map (
            O => \N__1136\,
            I => \un1_rData_0_sqmuxa_0\
        );

    \I__155\ : LocalMux
    port map (
            O => \N__1133\,
            I => \un1_rData_0_sqmuxa_0\
        );

    \I__154\ : InMux
    port map (
            O => \N__1128\,
            I => \N__1122\
        );

    \I__153\ : InMux
    port map (
            O => \N__1127\,
            I => \N__1122\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1122\,
            I => \rDataCounter_0_sqmuxa\
        );

    \I__151\ : IoInMux
    port map (
            O => \N__1119\,
            I => \N__1116\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1116\,
            I => \N__1113\
        );

    \I__149\ : IoSpan4Mux
    port map (
            O => \N__1113\,
            I => \N__1110\
        );

    \I__148\ : Span4Mux_s1_h
    port map (
            O => \N__1110\,
            I => \N__1107\
        );

    \I__147\ : Span4Mux_v
    port map (
            O => \N__1107\,
            I => \N__1104\
        );

    \I__146\ : Odrv4
    port map (
            O => \N__1104\,
            I => \oData_c_4\
        );

    \I__145\ : CascadeMux
    port map (
            O => \N__1101\,
            I => \rDatace_1_4_cascade_\
        );

    \I__144\ : CEMux
    port map (
            O => \N__1098\,
            I => \N__1095\
        );

    \I__143\ : LocalMux
    port map (
            O => \N__1095\,
            I => \rData_RNOZ0Z_4\
        );

    \I__142\ : CascadeMux
    port map (
            O => \N__1092\,
            I => \rDatace_1_5_cascade_\
        );

    \I__141\ : CEMux
    port map (
            O => \N__1089\,
            I => \N__1086\
        );

    \I__140\ : LocalMux
    port map (
            O => \N__1086\,
            I => \N__1083\
        );

    \I__139\ : Span4Mux_v
    port map (
            O => \N__1083\,
            I => \N__1080\
        );

    \I__138\ : Span4Mux_s1_h
    port map (
            O => \N__1080\,
            I => \N__1077\
        );

    \I__137\ : Odrv4
    port map (
            O => \N__1077\,
            I => \rData_RNOZ0Z_5\
        );

    \I__136\ : IoInMux
    port map (
            O => \N__1074\,
            I => \N__1071\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__1071\,
            I => \oData_c_2\
        );

    \I__134\ : CascadeMux
    port map (
            O => \N__1068\,
            I => \rDatace_1_0_cascade_\
        );

    \I__133\ : CEMux
    port map (
            O => \N__1065\,
            I => \N__1062\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__1062\,
            I => \rData_RNOZ0Z_0\
        );

    \I__131\ : CascadeMux
    port map (
            O => \N__1059\,
            I => \rDatace_1_1_cascade_\
        );

    \I__130\ : CEMux
    port map (
            O => \N__1056\,
            I => \N__1053\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__1053\,
            I => \N__1050\
        );

    \I__128\ : Span4Mux_s2_h
    port map (
            O => \N__1050\,
            I => \N__1047\
        );

    \I__127\ : Odrv4
    port map (
            O => \N__1047\,
            I => \rData_RNOZ0Z_1\
        );

    \I__126\ : CascadeMux
    port map (
            O => \N__1044\,
            I => \rDataCounter_0_sqmuxa_cascade_\
        );

    \I__125\ : CascadeMux
    port map (
            O => \N__1041\,
            I => \rDataCounter_RNO_0Z0Z_2_cascade_\
        );

    \I__124\ : InMux
    port map (
            O => \N__1038\,
            I => \rCycleCounter_cry_0\
        );

    \I__123\ : InMux
    port map (
            O => \N__1035\,
            I => \N__1032\
        );

    \I__122\ : LocalMux
    port map (
            O => \N__1032\,
            I => \rCycleCounter_s_2\
        );

    \I__121\ : InMux
    port map (
            O => \N__1029\,
            I => \rCycleCounter_cry_1\
        );

    \I__120\ : InMux
    port map (
            O => \N__1026\,
            I => \N__1023\
        );

    \I__119\ : LocalMux
    port map (
            O => \N__1023\,
            I => \N__1020\
        );

    \I__118\ : Odrv4
    port map (
            O => \N__1020\,
            I => \rCycleCounter_s_3\
        );

    \I__117\ : InMux
    port map (
            O => \N__1017\,
            I => \rCycleCounter_cry_2\
        );

    \I__116\ : CascadeMux
    port map (
            O => \N__1014\,
            I => \N__1010\
        );

    \I__115\ : InMux
    port map (
            O => \N__1013\,
            I => \N__1006\
        );

    \I__114\ : InMux
    port map (
            O => \N__1010\,
            I => \N__1001\
        );

    \I__113\ : InMux
    port map (
            O => \N__1009\,
            I => \N__1001\
        );

    \I__112\ : LocalMux
    port map (
            O => \N__1006\,
            I => \rCycleCounterZ0Z_4\
        );

    \I__111\ : LocalMux
    port map (
            O => \N__1001\,
            I => \rCycleCounterZ0Z_4\
        );

    \I__110\ : InMux
    port map (
            O => \N__996\,
            I => \N__993\
        );

    \I__109\ : LocalMux
    port map (
            O => \N__993\,
            I => \rCycleCounter_cry_3_THRU_CO\
        );

    \I__108\ : InMux
    port map (
            O => \N__990\,
            I => \rCycleCounter_cry_3\
        );

    \I__107\ : CascadeMux
    port map (
            O => \N__987\,
            I => \N__983\
        );

    \I__106\ : InMux
    port map (
            O => \N__986\,
            I => \N__980\
        );

    \I__105\ : InMux
    port map (
            O => \N__983\,
            I => \N__977\
        );

    \I__104\ : LocalMux
    port map (
            O => \N__980\,
            I => \rCycleCounterZ0Z_5\
        );

    \I__103\ : LocalMux
    port map (
            O => \N__977\,
            I => \rCycleCounterZ0Z_5\
        );

    \I__102\ : InMux
    port map (
            O => \N__972\,
            I => \N__969\
        );

    \I__101\ : LocalMux
    port map (
            O => \N__969\,
            I => \rCycleCounter_s_5\
        );

    \I__100\ : InMux
    port map (
            O => \N__966\,
            I => \rCycleCounter_cry_4\
        );

    \I__99\ : InMux
    port map (
            O => \N__963\,
            I => \N__959\
        );

    \I__98\ : InMux
    port map (
            O => \N__962\,
            I => \N__956\
        );

    \I__97\ : LocalMux
    port map (
            O => \N__959\,
            I => \rCycleCounterZ0Z_6\
        );

    \I__96\ : LocalMux
    port map (
            O => \N__956\,
            I => \rCycleCounterZ0Z_6\
        );

    \I__95\ : InMux
    port map (
            O => \N__951\,
            I => \N__948\
        );

    \I__94\ : LocalMux
    port map (
            O => \N__948\,
            I => \rCycleCounter_s_6\
        );

    \I__93\ : InMux
    port map (
            O => \N__945\,
            I => \rCycleCounter_cry_5\
        );

    \I__92\ : InMux
    port map (
            O => \N__942\,
            I => \rCycleCounter_cry_6\
        );

    \I__91\ : CascadeMux
    port map (
            O => \N__939\,
            I => \N__936\
        );

    \I__90\ : InMux
    port map (
            O => \N__936\,
            I => \N__932\
        );

    \I__89\ : InMux
    port map (
            O => \N__935\,
            I => \N__929\
        );

    \I__88\ : LocalMux
    port map (
            O => \N__932\,
            I => \rCycleCounterZ0Z_7\
        );

    \I__87\ : LocalMux
    port map (
            O => \N__929\,
            I => \rCycleCounterZ0Z_7\
        );

    \I__86\ : IoInMux
    port map (
            O => \N__924\,
            I => \N__921\
        );

    \I__85\ : LocalMux
    port map (
            O => \N__921\,
            I => \N__918\
        );

    \I__84\ : Odrv12
    port map (
            O => \N__918\,
            I => \oData_c_5\
        );

    \I__83\ : IoInMux
    port map (
            O => \N__915\,
            I => \N__912\
        );

    \I__82\ : LocalMux
    port map (
            O => \N__912\,
            I => \oData_c_1\
        );

    \I__81\ : CascadeMux
    port map (
            O => \N__909\,
            I => \pReceive_un12_rstate_3_cascade_\
        );

    \I__80\ : CascadeMux
    port map (
            O => \N__906\,
            I => \N_97_0_i_0_cascade_\
        );

    \I__79\ : IoInMux
    port map (
            O => \N__903\,
            I => \N__900\
        );

    \I__78\ : LocalMux
    port map (
            O => \N__900\,
            I => \oData_c_0\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \rData_0_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1898\,
            lcout => \oData_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1820\,
            ce => \N__1065\,
            sr => \_gnd_net_\
        );

    \rData_1_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1933\,
            lcout => \oData_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1818\,
            ce => \N__1056\,
            sr => \_gnd_net_\
        );

    \rCycleCounter_6_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110001100"
        )
    port map (
            in0 => \N__2085\,
            in1 => \N__1758\,
            in2 => \N__1969\,
            in3 => \N__951\,
            lcout => \rCycleCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1819\,
            ce => \N__1652\,
            sr => \_gnd_net_\
        );

    \rCycleCounter_4_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000111101011"
        )
    port map (
            in0 => \N__1759\,
            in1 => \N__996\,
            in2 => \N__1014\,
            in3 => \N__1140\,
            lcout => \rCycleCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1819\,
            ce => \N__1652\,
            sr => \_gnd_net_\
        );

    \rCycleCounter_5_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__1691\,
            in1 => \N__972\,
            in2 => \N__1968\,
            in3 => \N__1757\,
            lcout => \rCycleCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1819\,
            ce => \N__1652\,
            sr => \_gnd_net_\
        );

    \rCycleCounter_RNIPHLR_2_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1175\,
            in2 => \_gnd_net_\,
            in3 => \N__1199\,
            lcout => OPEN,
            ltout => \pReceive_un12_rstate_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_fast_RNIEUBD4_0_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__1689\,
            in1 => \N__1242\,
            in2 => \N__909\,
            in3 => \N__1155\,
            lcout => \N_97_0_i_0\,
            ltout => \N_97_0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_2_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__1934\,
            in1 => \N__1035\,
            in2 => \N__906\,
            in3 => \N__1690\,
            lcout => \rCycleCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1819\,
            ce => \N__1652\,
            sr => \_gnd_net_\
        );

    \rCycleCounter_3_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111001100"
        )
    port map (
            in0 => \N__2084\,
            in1 => \N__1026\,
            in2 => \N__1967\,
            in3 => \N__1756\,
            lcout => \rCycleCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1819\,
            ce => \N__1652\,
            sr => \_gnd_net_\
        );

    \rCycleCounter_RNIUFBN1_7_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1009\,
            in1 => \N__935\,
            in2 => \N__987\,
            in3 => \N__962\,
            lcout => \pReceive_un12_rstate_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_cry_c_0_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1233\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \rCycleCounter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_cry_0_THRU_LUT4_0_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1722\,
            in2 => \N__1308\,
            in3 => \N__1038\,
            lcout => \rCycleCounter_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \rCycleCounter_cry_0\,
            carryout => \rCycleCounter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_RNO_0_2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1198\,
            in2 => \N__1304\,
            in3 => \N__1029\,
            lcout => \rCycleCounter_s_2\,
            ltout => OPEN,
            carryin => \rCycleCounter_cry_1\,
            carryout => \rCycleCounter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_RNO_0_3_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1291\,
            in2 => \N__1179\,
            in3 => \N__1017\,
            lcout => \rCycleCounter_s_3\,
            ltout => OPEN,
            carryin => \rCycleCounter_cry_2\,
            carryout => \rCycleCounter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_cry_3_THRU_LUT4_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1013\,
            in2 => \N__1306\,
            in3 => \N__990\,
            lcout => \rCycleCounter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \rCycleCounter_cry_3\,
            carryout => \rCycleCounter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_RNO_0_5_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__986\,
            in2 => \N__1307\,
            in3 => \N__966\,
            lcout => \rCycleCounter_s_5\,
            ltout => OPEN,
            carryin => \rCycleCounter_cry_4\,
            carryout => \rCycleCounter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_RNO_0_6_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__963\,
            in2 => \N__1305\,
            in3 => \N__945\,
            lcout => \rCycleCounter_s_6\,
            ltout => OPEN,
            carryin => \rCycleCounter_cry_5\,
            carryout => \rCycleCounter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_7_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000100111"
        )
    port map (
            in0 => \N__1760\,
            in1 => \N__1139\,
            in2 => \N__939\,
            in3 => \N__942\,
            lcout => \rCycleCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1821\,
            ce => \N__1653\,
            sr => \_gnd_net_\
        );

    \rData_5_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1944\,
            lcout => \oData_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1824\,
            ce => \N__1089\,
            sr => \_gnd_net_\
        );

    \rData_2_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__1966\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \oData_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1827\,
            ce => \N__1254\,
            sr => \_gnd_net_\
        );

    \rData_RNO_0_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__1557\,
            in1 => \N__1502\,
            in2 => \_gnd_net_\,
            in3 => \N__1449\,
            lcout => OPEN,
            ltout => \rDatace_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_0_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__1389\,
            in1 => \N__1612\,
            in2 => \N__1068\,
            in3 => \N__2227\,
            lcout => \rData_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_0_1_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__1558\,
            in1 => \N__1503\,
            in2 => \_gnd_net_\,
            in3 => \N__1448\,
            lcout => OPEN,
            ltout => \rDatace_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__1390\,
            in1 => \N__1611\,
            in2 => \N__1059\,
            in3 => \N__2226\,
            lcout => \rData_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_0_2_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__1556\,
            in1 => \N__1501\,
            in2 => \_gnd_net_\,
            in3 => \N__1447\,
            lcout => \rDatace_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_0_rep1_RNIU3065_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__1619\,
            in1 => \N__2252\,
            in2 => \N__1406\,
            in3 => \N__2228\,
            lcout => \rDataCounter_0_sqmuxa\,
            ltout => \rDataCounter_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rDataCounter_1_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111111000"
        )
    port map (
            in0 => \N__2231\,
            in1 => \N__1668\,
            in2 => \N__1044\,
            in3 => \N__1508\,
            lcout => \rDataCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1822\,
            ce => 'H',
            sr => \N__1695\
        );

    \rDataCounter_RNO_0_2_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__1507\,
            in1 => \N__1667\,
            in2 => \N__1562\,
            in3 => \N__2229\,
            lcout => OPEN,
            ltout => \rDataCounter_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rDataCounter_2_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1041\,
            in3 => \N__1127\,
            lcout => \rDataCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1822\,
            ce => 'H',
            sr => \N__1695\
        );

    \rCycleCounter_RNIEVAN1_0_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1718\,
            in1 => \N__1226\,
            in2 => \N__1203\,
            in3 => \N__1174\,
            lcout => OPEN,
            ltout => \rCycleCounter_RNIEVAN1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_RNICFME3_0_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1158\,
            in3 => \N__1154\,
            lcout => \N_97_0_i\,
            ltout => \N_97_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_0_rep1_RNIDT874_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110011101"
        )
    port map (
            in0 => \N__1620\,
            in1 => \N__1398\,
            in2 => \N__1143\,
            in3 => \N__1927\,
            lcout => \un1_rData_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rDataCounter_0_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111010010"
        )
    port map (
            in0 => \N__2230\,
            in1 => \N__2169\,
            in2 => \N__1463\,
            in3 => \N__1128\,
            lcout => \rDataCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1822\,
            ce => 'H',
            sr => \N__1695\
        );

    \rData_4_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__1928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \oData_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1825\,
            ce => \N__1098\,
            sr => \_gnd_net_\
        );

    \rData_RNO_0_4_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__1540\,
            in1 => \N__1498\,
            in2 => \_gnd_net_\,
            in3 => \N__1446\,
            lcout => OPEN,
            ltout => \rDatace_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_4_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2161\,
            in1 => \N__1402\,
            in2 => \N__1101\,
            in3 => \N__2225\,
            lcout => \rData_RNOZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_0_5_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__1541\,
            in1 => \N__1499\,
            in2 => \_gnd_net_\,
            in3 => \N__1444\,
            lcout => OPEN,
            ltout => \rDatace_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_5_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2162\,
            in1 => \N__2072\,
            in2 => \N__1092\,
            in3 => \N__2223\,
            lcout => \rData_RNOZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_0_6_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__1542\,
            in1 => \N__1500\,
            in2 => \_gnd_net_\,
            in3 => \N__1445\,
            lcout => OPEN,
            ltout => \rDatace_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_6_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2163\,
            in1 => \N__2073\,
            in2 => \N__1332\,
            in3 => \N__2224\,
            lcout => \rData_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rDataCounter_RNIVRLB1_2_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__1539\,
            in1 => \N__1497\,
            in2 => \_gnd_net_\,
            in3 => \N__1443\,
            lcout => \pReceive_rdata_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_6_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1932\,
            lcout => \oData_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1828\,
            ce => \N__1317\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_2_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__1263\,
            in1 => \N__1613\,
            in2 => \N__1407\,
            in3 => \N__2239\,
            lcout => \rData_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_1_rep1_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__1970\,
            in1 => \N__2167\,
            in2 => \_gnd_net_\,
            in3 => \N__1382\,
            lcout => \rState_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1823\,
            ce => \N__2007\,
            sr => \_gnd_net_\
        );

    \rState_fast_RNI650B1_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__2021\,
            in1 => \N__1716\,
            in2 => \N__2103\,
            in3 => \N__1224\,
            lcout => g0_sn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rCycleCounter_0_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__1225\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1766\,
            lcout => \rCycleCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1829\,
            ce => \N__1634\,
            sr => \_gnd_net_\
        );

    \rCycleCounter_1_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__1767\,
            in1 => \N__1734\,
            in2 => \_gnd_net_\,
            in3 => \N__1717\,
            lcout => \rCycleCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1829\,
            ce => \N__1634\,
            sr => \_gnd_net_\
        );

    \rState_fast_RNIHNAF_0_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2101\,
            in2 => \_gnd_net_\,
            in3 => \N__2020\,
            lcout => \pReceive_rstate\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_0_rep1_RNIDN6N_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__1595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1462\,
            lcout => \CO0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_0_rep1_RNIJOJB_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1594\,
            in2 => \_gnd_net_\,
            in3 => \N__1368\,
            lcout => \rCycleCountere_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_0_rep1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__1599\,
            in1 => \N__2066\,
            in2 => \_gnd_net_\,
            in3 => \N__1974\,
            lcout => \rState_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1830\,
            ce => \N__2006\,
            sr => \_gnd_net_\
        );

    \rState_0_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101111"
        )
    port map (
            in0 => \N__2067\,
            in1 => \_gnd_net_\,
            in2 => \N__1986\,
            in3 => \N__2153\,
            lcout => \rStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1830\,
            ce => \N__2006\,
            sr => \_gnd_net_\
        );

    \rState_1_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010110101010"
        )
    port map (
            in0 => \N__2068\,
            in1 => \_gnd_net_\,
            in2 => \N__1987\,
            in3 => \N__2154\,
            lcout => \rStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1830\,
            ce => \N__2006\,
            sr => \_gnd_net_\
        );

    \rData_RNO_0_3_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__1563\,
            in1 => \N__1512\,
            in2 => \_gnd_net_\,
            in3 => \N__1464\,
            lcout => OPEN,
            ltout => \rDatace_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_3_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2139\,
            in1 => \N__1397\,
            in2 => \N__1335\,
            in3 => \N__2241\,
            lcout => \rData_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_3_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1988\,
            lcout => \oData_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1833\,
            ce => \N__2292\,
            sr => \_gnd_net_\
        );

    \rDataReady_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__2273\,
            in1 => \N__2078\,
            in2 => \_gnd_net_\,
            in3 => \N__2168\,
            lcout => \oDataReady_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_RNI2GHJ5_1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010110011"
        )
    port map (
            in0 => \N__2262\,
            in1 => \N__2064\,
            in2 => \N__2240\,
            in3 => \N__2151\,
            lcout => \un1_rCycleCounter_2_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rData_RNO_7_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2150\,
            in1 => \N__2261\,
            in2 => \N__2077\,
            in3 => \N__2232\,
            lcout => \rData_RNOZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rState_fast_1_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011000100110"
        )
    port map (
            in0 => \N__2102\,
            in1 => \N__2152\,
            in2 => \N__1989\,
            in3 => \_gnd_net_\,
            lcout => \rState_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1831\,
            ce => \N__2005\,
            sr => \_gnd_net_\
        );

    \rState_fast_0_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__2065\,
            in1 => \N__1982\,
            in2 => \_gnd_net_\,
            in3 => \N__2022\,
            lcout => \rState_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1831\,
            ce => \N__2005\,
            sr => \_gnd_net_\
        );

    \rData_7_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__1978\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \oData_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1832\,
            ce => \N__1779\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
